//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Sat Sep 09 16:40:21 2023

module Gowin_SDPB (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [5:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [16:0] ada;
input [5:0] din;
input [16:0] adb;

wire lut_f_0;
wire lut_f_1;
wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [0:0] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [0:0] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [0:0] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [1:1] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [1:1] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [1:1] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [1:1] sdpb_inst_7_dout;
wire [30:0] sdpb_inst_8_dout_w;
wire [2:2] sdpb_inst_8_dout;
wire [30:0] sdpb_inst_9_dout_w;
wire [2:2] sdpb_inst_9_dout;
wire [30:0] sdpb_inst_10_dout_w;
wire [2:2] sdpb_inst_10_dout;
wire [30:0] sdpb_inst_11_dout_w;
wire [2:2] sdpb_inst_11_dout;
wire [30:0] sdpb_inst_12_dout_w;
wire [3:3] sdpb_inst_12_dout;
wire [30:0] sdpb_inst_13_dout_w;
wire [3:3] sdpb_inst_13_dout;
wire [30:0] sdpb_inst_14_dout_w;
wire [3:3] sdpb_inst_14_dout;
wire [30:0] sdpb_inst_15_dout_w;
wire [3:3] sdpb_inst_15_dout;
wire [30:0] sdpb_inst_16_dout_w;
wire [4:4] sdpb_inst_16_dout;
wire [30:0] sdpb_inst_17_dout_w;
wire [4:4] sdpb_inst_17_dout;
wire [30:0] sdpb_inst_18_dout_w;
wire [4:4] sdpb_inst_18_dout;
wire [30:0] sdpb_inst_19_dout_w;
wire [4:4] sdpb_inst_19_dout;
wire [30:0] sdpb_inst_20_dout_w;
wire [5:5] sdpb_inst_20_dout;
wire [30:0] sdpb_inst_21_dout_w;
wire [5:5] sdpb_inst_21_dout;
wire [30:0] sdpb_inst_22_dout_w;
wire [5:5] sdpb_inst_22_dout;
wire [30:0] sdpb_inst_23_dout_w;
wire [5:5] sdpb_inst_23_dout;
wire [30:0] sdpb_inst_24_dout_w;
wire [0:0] sdpb_inst_24_dout;
wire [30:0] sdpb_inst_25_dout_w;
wire [0:0] sdpb_inst_25_dout;
wire [30:0] sdpb_inst_26_dout_w;
wire [1:1] sdpb_inst_26_dout;
wire [30:0] sdpb_inst_27_dout_w;
wire [1:1] sdpb_inst_27_dout;
wire [30:0] sdpb_inst_28_dout_w;
wire [2:2] sdpb_inst_28_dout;
wire [30:0] sdpb_inst_29_dout_w;
wire [2:2] sdpb_inst_29_dout;
wire [30:0] sdpb_inst_30_dout_w;
wire [3:3] sdpb_inst_30_dout;
wire [30:0] sdpb_inst_31_dout_w;
wire [3:3] sdpb_inst_31_dout;
wire [30:0] sdpb_inst_32_dout_w;
wire [4:4] sdpb_inst_32_dout;
wire [30:0] sdpb_inst_33_dout_w;
wire [4:4] sdpb_inst_33_dout;
wire [30:0] sdpb_inst_34_dout_w;
wire [5:5] sdpb_inst_34_dout;
wire [30:0] sdpb_inst_35_dout_w;
wire [5:5] sdpb_inst_35_dout;
wire [30:0] sdpb_inst_36_dout_w;
wire [0:0] sdpb_inst_36_dout;
wire [30:0] sdpb_inst_37_dout_w;
wire [1:1] sdpb_inst_37_dout;
wire [30:0] sdpb_inst_38_dout_w;
wire [2:2] sdpb_inst_38_dout;
wire [30:0] sdpb_inst_39_dout_w;
wire [3:3] sdpb_inst_39_dout;
wire [30:0] sdpb_inst_40_dout_w;
wire [4:4] sdpb_inst_40_dout;
wire [30:0] sdpb_inst_41_dout_w;
wire [5:5] sdpb_inst_41_dout;
wire [25:0] sdpb_inst_42_dout_w;
wire [5:0] sdpb_inst_42_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT6 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14]),
  .I4(ada[15]),
  .I5(ada[16])
);
defparam lut_inst_0.INIT = 64'h0100000000000000;
LUT6 lut_inst_1 (
  .F(lut_f_1),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14]),
  .I4(adb[15]),
  .I5(adb[16])
);
defparam lut_inst_1.INIT = 64'h0100000000000000;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_2.RESET_MODE = "SYNC";

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_3.RESET_MODE = "SYNC";

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_4.RESET_MODE = "SYNC";

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b0;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_5.RESET_MODE = "SYNC";

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b0;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_6.RESET_MODE = "SYNC";

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b0;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_7.RESET_MODE = "SYNC";

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[30:0],sdpb_inst_8_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_8.READ_MODE = 1'b0;
defparam sdpb_inst_8.BIT_WIDTH_0 = 1;
defparam sdpb_inst_8.BIT_WIDTH_1 = 1;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_8.RESET_MODE = "SYNC";

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[30:0],sdpb_inst_9_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_9.READ_MODE = 1'b0;
defparam sdpb_inst_9.BIT_WIDTH_0 = 1;
defparam sdpb_inst_9.BIT_WIDTH_1 = 1;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_9.RESET_MODE = "SYNC";

SDPB sdpb_inst_10 (
    .DO({sdpb_inst_10_dout_w[30:0],sdpb_inst_10_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_10.READ_MODE = 1'b0;
defparam sdpb_inst_10.BIT_WIDTH_0 = 1;
defparam sdpb_inst_10.BIT_WIDTH_1 = 1;
defparam sdpb_inst_10.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_10.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_10.RESET_MODE = "SYNC";

SDPB sdpb_inst_11 (
    .DO({sdpb_inst_11_dout_w[30:0],sdpb_inst_11_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_11.READ_MODE = 1'b0;
defparam sdpb_inst_11.BIT_WIDTH_0 = 1;
defparam sdpb_inst_11.BIT_WIDTH_1 = 1;
defparam sdpb_inst_11.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_11.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_11.RESET_MODE = "SYNC";

SDPB sdpb_inst_12 (
    .DO({sdpb_inst_12_dout_w[30:0],sdpb_inst_12_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_12.READ_MODE = 1'b0;
defparam sdpb_inst_12.BIT_WIDTH_0 = 1;
defparam sdpb_inst_12.BIT_WIDTH_1 = 1;
defparam sdpb_inst_12.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_12.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_12.RESET_MODE = "SYNC";

SDPB sdpb_inst_13 (
    .DO({sdpb_inst_13_dout_w[30:0],sdpb_inst_13_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_13.READ_MODE = 1'b0;
defparam sdpb_inst_13.BIT_WIDTH_0 = 1;
defparam sdpb_inst_13.BIT_WIDTH_1 = 1;
defparam sdpb_inst_13.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_13.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_13.RESET_MODE = "SYNC";

SDPB sdpb_inst_14 (
    .DO({sdpb_inst_14_dout_w[30:0],sdpb_inst_14_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_14.READ_MODE = 1'b0;
defparam sdpb_inst_14.BIT_WIDTH_0 = 1;
defparam sdpb_inst_14.BIT_WIDTH_1 = 1;
defparam sdpb_inst_14.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_14.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_14.RESET_MODE = "SYNC";

SDPB sdpb_inst_15 (
    .DO({sdpb_inst_15_dout_w[30:0],sdpb_inst_15_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_15.READ_MODE = 1'b0;
defparam sdpb_inst_15.BIT_WIDTH_0 = 1;
defparam sdpb_inst_15.BIT_WIDTH_1 = 1;
defparam sdpb_inst_15.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_15.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_15.RESET_MODE = "SYNC";

SDPB sdpb_inst_16 (
    .DO({sdpb_inst_16_dout_w[30:0],sdpb_inst_16_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_16.READ_MODE = 1'b0;
defparam sdpb_inst_16.BIT_WIDTH_0 = 1;
defparam sdpb_inst_16.BIT_WIDTH_1 = 1;
defparam sdpb_inst_16.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_16.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_16.RESET_MODE = "SYNC";

SDPB sdpb_inst_17 (
    .DO({sdpb_inst_17_dout_w[30:0],sdpb_inst_17_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_17.READ_MODE = 1'b0;
defparam sdpb_inst_17.BIT_WIDTH_0 = 1;
defparam sdpb_inst_17.BIT_WIDTH_1 = 1;
defparam sdpb_inst_17.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_17.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_17.RESET_MODE = "SYNC";

SDPB sdpb_inst_18 (
    .DO({sdpb_inst_18_dout_w[30:0],sdpb_inst_18_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_18.READ_MODE = 1'b0;
defparam sdpb_inst_18.BIT_WIDTH_0 = 1;
defparam sdpb_inst_18.BIT_WIDTH_1 = 1;
defparam sdpb_inst_18.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_18.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_18.RESET_MODE = "SYNC";

SDPB sdpb_inst_19 (
    .DO({sdpb_inst_19_dout_w[30:0],sdpb_inst_19_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_19.READ_MODE = 1'b0;
defparam sdpb_inst_19.BIT_WIDTH_0 = 1;
defparam sdpb_inst_19.BIT_WIDTH_1 = 1;
defparam sdpb_inst_19.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_19.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_19.RESET_MODE = "SYNC";

SDPB sdpb_inst_20 (
    .DO({sdpb_inst_20_dout_w[30:0],sdpb_inst_20_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_20.READ_MODE = 1'b0;
defparam sdpb_inst_20.BIT_WIDTH_0 = 1;
defparam sdpb_inst_20.BIT_WIDTH_1 = 1;
defparam sdpb_inst_20.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_20.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_20.RESET_MODE = "SYNC";

SDPB sdpb_inst_21 (
    .DO({sdpb_inst_21_dout_w[30:0],sdpb_inst_21_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_21.READ_MODE = 1'b0;
defparam sdpb_inst_21.BIT_WIDTH_0 = 1;
defparam sdpb_inst_21.BIT_WIDTH_1 = 1;
defparam sdpb_inst_21.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_21.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_21.RESET_MODE = "SYNC";

SDPB sdpb_inst_22 (
    .DO({sdpb_inst_22_dout_w[30:0],sdpb_inst_22_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_22.READ_MODE = 1'b0;
defparam sdpb_inst_22.BIT_WIDTH_0 = 1;
defparam sdpb_inst_22.BIT_WIDTH_1 = 1;
defparam sdpb_inst_22.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_22.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_22.RESET_MODE = "SYNC";

SDPB sdpb_inst_23 (
    .DO({sdpb_inst_23_dout_w[30:0],sdpb_inst_23_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_23.READ_MODE = 1'b0;
defparam sdpb_inst_23.BIT_WIDTH_0 = 1;
defparam sdpb_inst_23.BIT_WIDTH_1 = 1;
defparam sdpb_inst_23.BLK_SEL_0 = 3'b011;
defparam sdpb_inst_23.BLK_SEL_1 = 3'b011;
defparam sdpb_inst_23.RESET_MODE = "SYNC";

SDPB sdpb_inst_24 (
    .DO({sdpb_inst_24_dout_w[30:0],sdpb_inst_24_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_24.READ_MODE = 1'b0;
defparam sdpb_inst_24.BIT_WIDTH_0 = 1;
defparam sdpb_inst_24.BIT_WIDTH_1 = 1;
defparam sdpb_inst_24.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_24.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_24.RESET_MODE = "SYNC";

SDPB sdpb_inst_25 (
    .DO({sdpb_inst_25_dout_w[30:0],sdpb_inst_25_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_25.READ_MODE = 1'b0;
defparam sdpb_inst_25.BIT_WIDTH_0 = 1;
defparam sdpb_inst_25.BIT_WIDTH_1 = 1;
defparam sdpb_inst_25.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_25.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_25.RESET_MODE = "SYNC";

SDPB sdpb_inst_26 (
    .DO({sdpb_inst_26_dout_w[30:0],sdpb_inst_26_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_26.READ_MODE = 1'b0;
defparam sdpb_inst_26.BIT_WIDTH_0 = 1;
defparam sdpb_inst_26.BIT_WIDTH_1 = 1;
defparam sdpb_inst_26.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_26.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_26.RESET_MODE = "SYNC";

SDPB sdpb_inst_27 (
    .DO({sdpb_inst_27_dout_w[30:0],sdpb_inst_27_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_27.READ_MODE = 1'b0;
defparam sdpb_inst_27.BIT_WIDTH_0 = 1;
defparam sdpb_inst_27.BIT_WIDTH_1 = 1;
defparam sdpb_inst_27.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_27.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_27.RESET_MODE = "SYNC";

SDPB sdpb_inst_28 (
    .DO({sdpb_inst_28_dout_w[30:0],sdpb_inst_28_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_28.READ_MODE = 1'b0;
defparam sdpb_inst_28.BIT_WIDTH_0 = 1;
defparam sdpb_inst_28.BIT_WIDTH_1 = 1;
defparam sdpb_inst_28.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_28.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_28.RESET_MODE = "SYNC";

SDPB sdpb_inst_29 (
    .DO({sdpb_inst_29_dout_w[30:0],sdpb_inst_29_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_29.READ_MODE = 1'b0;
defparam sdpb_inst_29.BIT_WIDTH_0 = 1;
defparam sdpb_inst_29.BIT_WIDTH_1 = 1;
defparam sdpb_inst_29.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_29.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_29.RESET_MODE = "SYNC";

SDPB sdpb_inst_30 (
    .DO({sdpb_inst_30_dout_w[30:0],sdpb_inst_30_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_30.READ_MODE = 1'b0;
defparam sdpb_inst_30.BIT_WIDTH_0 = 1;
defparam sdpb_inst_30.BIT_WIDTH_1 = 1;
defparam sdpb_inst_30.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_30.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_30.RESET_MODE = "SYNC";

SDPB sdpb_inst_31 (
    .DO({sdpb_inst_31_dout_w[30:0],sdpb_inst_31_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_31.READ_MODE = 1'b0;
defparam sdpb_inst_31.BIT_WIDTH_0 = 1;
defparam sdpb_inst_31.BIT_WIDTH_1 = 1;
defparam sdpb_inst_31.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_31.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_31.RESET_MODE = "SYNC";

SDPB sdpb_inst_32 (
    .DO({sdpb_inst_32_dout_w[30:0],sdpb_inst_32_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_32.READ_MODE = 1'b0;
defparam sdpb_inst_32.BIT_WIDTH_0 = 1;
defparam sdpb_inst_32.BIT_WIDTH_1 = 1;
defparam sdpb_inst_32.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_32.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_32.RESET_MODE = "SYNC";

SDPB sdpb_inst_33 (
    .DO({sdpb_inst_33_dout_w[30:0],sdpb_inst_33_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_33.READ_MODE = 1'b0;
defparam sdpb_inst_33.BIT_WIDTH_0 = 1;
defparam sdpb_inst_33.BIT_WIDTH_1 = 1;
defparam sdpb_inst_33.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_33.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_33.RESET_MODE = "SYNC";

SDPB sdpb_inst_34 (
    .DO({sdpb_inst_34_dout_w[30:0],sdpb_inst_34_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_34.READ_MODE = 1'b0;
defparam sdpb_inst_34.BIT_WIDTH_0 = 1;
defparam sdpb_inst_34.BIT_WIDTH_1 = 1;
defparam sdpb_inst_34.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_34.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_34.RESET_MODE = "SYNC";

SDPB sdpb_inst_35 (
    .DO({sdpb_inst_35_dout_w[30:0],sdpb_inst_35_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_35.READ_MODE = 1'b0;
defparam sdpb_inst_35.BIT_WIDTH_0 = 1;
defparam sdpb_inst_35.BIT_WIDTH_1 = 1;
defparam sdpb_inst_35.BLK_SEL_0 = 3'b101;
defparam sdpb_inst_35.BLK_SEL_1 = 3'b101;
defparam sdpb_inst_35.RESET_MODE = "SYNC";

SDPB sdpb_inst_36 (
    .DO({sdpb_inst_36_dout_w[30:0],sdpb_inst_36_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_36.READ_MODE = 1'b0;
defparam sdpb_inst_36.BIT_WIDTH_0 = 1;
defparam sdpb_inst_36.BIT_WIDTH_1 = 1;
defparam sdpb_inst_36.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_36.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_36.RESET_MODE = "SYNC";

SDPB sdpb_inst_37 (
    .DO({sdpb_inst_37_dout_w[30:0],sdpb_inst_37_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_37.READ_MODE = 1'b0;
defparam sdpb_inst_37.BIT_WIDTH_0 = 1;
defparam sdpb_inst_37.BIT_WIDTH_1 = 1;
defparam sdpb_inst_37.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_37.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_37.RESET_MODE = "SYNC";

SDPB sdpb_inst_38 (
    .DO({sdpb_inst_38_dout_w[30:0],sdpb_inst_38_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_38.READ_MODE = 1'b0;
defparam sdpb_inst_38.BIT_WIDTH_0 = 1;
defparam sdpb_inst_38.BIT_WIDTH_1 = 1;
defparam sdpb_inst_38.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_38.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_38.RESET_MODE = "SYNC";

SDPB sdpb_inst_39 (
    .DO({sdpb_inst_39_dout_w[30:0],sdpb_inst_39_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_39.READ_MODE = 1'b0;
defparam sdpb_inst_39.BIT_WIDTH_0 = 1;
defparam sdpb_inst_39.BIT_WIDTH_1 = 1;
defparam sdpb_inst_39.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_39.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_39.RESET_MODE = "SYNC";

SDPB sdpb_inst_40 (
    .DO({sdpb_inst_40_dout_w[30:0],sdpb_inst_40_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_40.READ_MODE = 1'b0;
defparam sdpb_inst_40.BIT_WIDTH_0 = 1;
defparam sdpb_inst_40.BIT_WIDTH_1 = 1;
defparam sdpb_inst_40.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_40.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_40.RESET_MODE = "SYNC";

SDPB sdpb_inst_41 (
    .DO({sdpb_inst_41_dout_w[30:0],sdpb_inst_41_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[16],ada[15],ada[14]}),
    .BLKSELB({adb[16],adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_41.READ_MODE = 1'b0;
defparam sdpb_inst_41.BIT_WIDTH_0 = 1;
defparam sdpb_inst_41.BIT_WIDTH_1 = 1;
defparam sdpb_inst_41.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_41.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_41.RESET_MODE = "SYNC";

SDPB sdpb_inst_42 (
    .DO({sdpb_inst_42_dout_w[25:0],sdpb_inst_42_dout[5:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_1}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_42.READ_MODE = 1'b0;
defparam sdpb_inst_42.BIT_WIDTH_0 = 8;
defparam sdpb_inst_42.BIT_WIDTH_1 = 8;
defparam sdpb_inst_42.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_42.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_42.RESET_MODE = "SYNC";

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[16]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[15]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(sdpb_inst_2_dout[0]),
  .I1(sdpb_inst_3_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(sdpb_inst_24_dout[0]),
  .I1(sdpb_inst_25_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(sdpb_inst_36_dout[0]),
  .I1(sdpb_inst_42_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_24),
  .I1(mux_o_25),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(mux_o_26),
  .I1(mux_o_27),
  .S0(dff_q_1)
);
MUX2 mux_inst_30 (
  .O(dout[0]),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_0)
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(sdpb_inst_4_dout[1]),
  .I1(sdpb_inst_5_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(sdpb_inst_6_dout[1]),
  .I1(sdpb_inst_7_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(sdpb_inst_26_dout[1]),
  .I1(sdpb_inst_27_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(sdpb_inst_37_dout[1]),
  .I1(sdpb_inst_42_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(dff_q_1)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(dff_q_1)
);
MUX2 mux_inst_61 (
  .O(dout[1]),
  .I0(mux_o_59),
  .I1(mux_o_60),
  .S0(dff_q_0)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(sdpb_inst_8_dout[2]),
  .I1(sdpb_inst_9_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(sdpb_inst_10_dout[2]),
  .I1(sdpb_inst_11_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(sdpb_inst_28_dout[2]),
  .I1(sdpb_inst_29_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(sdpb_inst_38_dout[2]),
  .I1(sdpb_inst_42_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(dff_q_1)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(dff_q_1)
);
MUX2 mux_inst_92 (
  .O(dout[2]),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_0)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(sdpb_inst_12_dout[3]),
  .I1(sdpb_inst_13_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(sdpb_inst_14_dout[3]),
  .I1(sdpb_inst_15_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(sdpb_inst_30_dout[3]),
  .I1(sdpb_inst_31_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(sdpb_inst_39_dout[3]),
  .I1(sdpb_inst_42_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(dff_q_1)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(dff_q_1)
);
MUX2 mux_inst_123 (
  .O(dout[3]),
  .I0(mux_o_121),
  .I1(mux_o_122),
  .S0(dff_q_0)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(sdpb_inst_16_dout[4]),
  .I1(sdpb_inst_17_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(sdpb_inst_18_dout[4]),
  .I1(sdpb_inst_19_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(sdpb_inst_32_dout[4]),
  .I1(sdpb_inst_33_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(sdpb_inst_40_dout[4]),
  .I1(sdpb_inst_42_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(mux_o_148),
  .I1(mux_o_149),
  .S0(dff_q_1)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(dff_q_1)
);
MUX2 mux_inst_154 (
  .O(dout[4]),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(dff_q_0)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(sdpb_inst_20_dout[5]),
  .I1(sdpb_inst_21_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(sdpb_inst_22_dout[5]),
  .I1(sdpb_inst_23_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(sdpb_inst_34_dout[5]),
  .I1(sdpb_inst_35_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(sdpb_inst_41_dout[5]),
  .I1(sdpb_inst_42_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(dff_q_1)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_1)
);
MUX2 mux_inst_185 (
  .O(dout[5]),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(dff_q_0)
);
endmodule //Gowin_SDPB
