//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Thu Sep 07 10:46:34 2023

module Gowin_SDPB (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);//morhology_3x3v2

output [0:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [17:0] ada;
input [0:0] din;
input [17:0] adb;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [0:0] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [0:0] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [0:0] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [0:0] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [0:0] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [0:0] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [0:0] sdpb_inst_7_dout;
wire [30:0] sdpb_inst_8_dout_w;
wire [0:0] sdpb_inst_8_dout;
wire [30:0] sdpb_inst_9_dout_w;
wire [0:0] sdpb_inst_9_dout;
wire [30:0] sdpb_inst_10_dout_w;
wire [0:0] sdpb_inst_10_dout;
wire [30:0] sdpb_inst_11_dout_w;
wire [0:0] sdpb_inst_11_dout;
wire [30:0] sdpb_inst_12_dout_w;
wire [0:0] sdpb_inst_12_dout;
wire [30:0] sdpb_inst_13_dout_w;
wire [0:0] sdpb_inst_13_dout;
wire [30:0] sdpb_inst_14_dout_w;
wire [0:0] sdpb_inst_14_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire dff_q_7;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_8.INIT = 16'h0100;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_9.INIT = 16'h0200;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_10.INIT = 16'h0400;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_11.INIT = 16'h0800;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_12.INIT = 16'h1000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_13.INIT = 16'h2000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_14.INIT = 16'h4000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_15.INIT = 16'h0001;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_16.INIT = 16'h0002;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_17.INIT = 16'h0004;
LUT4 lut_inst_18 (
  .F(lut_f_18),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_18.INIT = 16'h0008;
LUT4 lut_inst_19 (
  .F(lut_f_19),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_19.INIT = 16'h0010;
LUT4 lut_inst_20 (
  .F(lut_f_20),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_20.INIT = 16'h0020;
LUT4 lut_inst_21 (
  .F(lut_f_21),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_21.INIT = 16'h0040;
LUT4 lut_inst_22 (
  .F(lut_f_22),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_22.INIT = 16'h0080;
LUT4 lut_inst_23 (
  .F(lut_f_23),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_23.INIT = 16'h0100;
LUT4 lut_inst_24 (
  .F(lut_f_24),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_24.INIT = 16'h0200;
LUT4 lut_inst_25 (
  .F(lut_f_25),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_25.INIT = 16'h0400;
LUT4 lut_inst_26 (
  .F(lut_f_26),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_26.INIT = 16'h0800;
LUT4 lut_inst_27 (
  .F(lut_f_27),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_27.INIT = 16'h1000;
LUT4 lut_inst_28 (
  .F(lut_f_28),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_28.INIT = 16'h2000;
LUT4 lut_inst_29 (
  .F(lut_f_29),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_29.INIT = 16'h4000;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_15}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b1;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_16}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b1;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFF;
defparam sdpb_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h9F0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1E = 256'hFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFCF803FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_20 = 256'hFFF818F83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFF807FF8FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_25 = 256'hFFFFFFF383FFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07FFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFE01FFFFFFFFFFFFFFFFFFFFFFF507FFFE3FFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2A = 256'hFFFFFFFFFFE70FFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007FFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFF001FFFFFFFFFFFFFFFFFFFFFFF9FFFFF0017FFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFF;
defparam sdpb_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFF400000FFF;
defparam sdpb_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFF;
defparam sdpb_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8400001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFC0007F;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_37 = 256'hF83FFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFF00000;
defparam sdpb_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h0007FFFFFFFFFFFFFFFFFFFFFFFFF000000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3C = 256'hFFFFFF803FFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sdpb_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3E = 256'hFFFBC0007FFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003FFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_17}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b1;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'hFFFE000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFF8F0001FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_03 = 256'hFFFFFFFC3C000FFFFFFFFFFFFFFFFFFFFFFFFF8000000007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_05 = 256'hFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFC0F0007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_08 = 256'hFFFFFFFFFFFE03C007FFFFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0A = 256'hFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFF00F003FFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFF003C03F3FFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFF;
defparam sdpb_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFF;
defparam sdpb_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8003E7FFFFFFFFFFFFFFFFF800F81F0FFFFFF;
defparam sdpb_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h0787FFFFFFFFFFFFFFFF8003E0F83FFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
defparam sdpb_inst_2.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam sdpb_inst_2.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001E07FFFFFFFFFFFFFFFC00078FC0F;
defparam sdpb_inst_2.INIT_RAM_16 = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_17 = 256'hFFFC007C07FFFFFFFFFFFFFFE0001F7C03FFFFFFFFFFFFFFFFFFFFFFFFFC0000;
defparam sdpb_inst_2.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_19 = 256'hFE00FFFFFFFFFFFFFFFFFFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00F007FFFFFFFFFFFFFF00007;
defparam sdpb_inst_2.INIT_RAM_1B = 256'hF00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1C = 256'hFFFFFFFFFC03C007FFFFFFFFFFFFFC0001FF003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h00007F000FFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFC0F8007FFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_20 = 256'hFFFFFFFC000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFF8FC1E0007FFFFFFFFFFFFC0001F8003FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_23 = 256'hFFF9F0000FC000FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FC78000FFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_25 = 256'hFFFFFFFFFFFFF8000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFC1F9F0001FFFFFFFFFFC3C0007F0003FFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_28 = 256'hFFFFFFFC0F8003F8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000FFFFFFF;
defparam sdpb_inst_2.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FFC0007FF;
defparam sdpb_inst_2.INIT_RAM_2A = 256'hFFFFFFFFF1FFFFFFFFE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFE01FF0001FFFFFFFFFE03E003FE0003FFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h007E7FFFFFFF00F801FF8000FFFFFFFFFFFFFFFFE1F01FFFFFFFFE000000003F;
defparam sdpb_inst_2.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF801FE0;
defparam sdpb_inst_2.INIT_RAM_2F = 256'hFFFFFFFFFFE0380383FFFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FC000F87FFFFFF003E00F9E0007FFFFF;
defparam sdpb_inst_2.INIT_RAM_31 = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_32 = 256'h003F8003E07FFFFF800F80FC78003FFFFFFFFFFFFFFFF00000807FFFFFF80000;
defparam sdpb_inst_2.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFC0000000FFFFFFF000000003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007F000F807FFFF8003E07E1E001F;
defparam sdpb_inst_2.INIT_RAM_36 = 256'hE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_37 = 256'hFFFFE000FF001F007FFFC000F83E07801FFFFFFFFFFFFFFF80000000030FFFFF;
defparam sdpb_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_39 = 256'hE00E3FFFFFFFFFFFFF800000000000FFFFFC000000007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FF007C007FFE0001FFF01;
defparam sdpb_inst_2.INIT_RAM_3B = 256'h1FFFFF8000000017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFF000F9F01F0007FE00007FF80780F0FFFFFFFFFFFFFE00000000000;
defparam sdpb_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3E = 256'hFF800E0783FFFFFFFFFFFFF0000000000007FFFFF000000004FFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001E1F03C0007F80001;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_18}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b1;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'h00000001FFFE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFC007C1F0F8000FC00007FC0038380FFFFFFFFFFFFFC0000F0;
defparam sdpb_inst_3.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_03 = 256'h80001FC000E1C03FFFFFFFFFFFF800007FFE0000003FFFC000000003FFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF801F03F3E0001F;
defparam sdpb_inst_3.INIT_RAM_05 = 256'h0FFFFFE000000FFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFF803C03EF80007E00007E0003DE00FFFFFFFFFFFFC00;
defparam sdpb_inst_3.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_08 = 256'h0000F80003F0000FF003FFFFFFFFFFFE0007FFFFFFE00001FFFF800000000FFF;
defparam sdpb_inst_3.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFF80F803FF;
defparam sdpb_inst_3.INIT_RAM_0A = 256'hFF8003FFFFFFFC00007FFFF000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0B = 256'hFFFFFFFFFFFFC00FFFFFFFFFFFF83E007FC0003E0001FC0003F000FFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0C = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0D = 256'h8007F8000F8000FF0000F8003FFFFFFFFFFFE003FFFFFFFFC00007FFFE000000;
defparam sdpb_inst_3.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFF001FFFFFFFFFF3F87;
defparam sdpb_inst_3.INIT_RAM_0F = 256'hFFFFFFF001FFFFFFFFFF80007FFFC100000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_10 = 256'hFFFFFFFFFFFE007FF8007FFFFFFFFFC3F9F0007F0003F000FFC0007C000FFFFF;
defparam sdpb_inst_3.INIT_RAM_11 = 256'h080000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_12 = 256'hF83FFC000FF000FC007FF0003F0003FFFFFFFFFFF8007FFFFFFFFFF0000FFFF8;
defparam sdpb_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FFE001FFE03FFFF;
defparam sdpb_inst_3.INIT_RAM_14 = 256'hFFFFFFFFFFFC003FFFFFFFFFFE0003FFFF060000000FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFC003FF8007FF007FFFFE03FF0003FE001F007E3E001FC001;
defparam sdpb_inst_3.INIT_RAM_16 = 256'h7FFFE040000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_17 = 256'h0FFFFFC03FE0007FE007C03E0F800FF000FFFFFFFFFFFE001FFFFFFFFFFFE000;
defparam sdpb_inst_3.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FFE000FFC0;
defparam sdpb_inst_3.INIT_RAM_19 = 256'hBC007FFFFFFFFFFF800FFFFFFFFFFFFE001FFFFC000000003FFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFC003FFC003FE003FFFFF003F8001EFE01F01F03E007;
defparam sdpb_inst_3.INIT_RAM_1B = 256'hFFC000FFFF8100000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1C = 256'h1FF800FFFFFC003F00079FE07E1F80F8078F003FFFFFFFFFFFE003FFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FF80;
defparam sdpb_inst_3.INIT_RAM_1E = 256'h3E03C3C01FFFFFFFFFFFF801FFFFFFFFFFFFF0000FFFF0000000007FFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFC3FC001FFF81FFE003FFFFF8007F000E1FE1F8F80;
defparam sdpb_inst_3.INIT_RAM_20 = 256'hFFFFFFFE0001FFFE000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_21 = 256'h7FFF87FF800FFFFFE001FF003C1FE3E7C00F81E0701FFFFFFFFFFFFE007FFFFF;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803FC00;
defparam sdpb_inst_3.INIT_RAM_23 = 256'hFFC003E1F01C0FFFFFFFFFFFFF803FFFFFFFFFFFFFC0007FFFC0000000018000;
defparam sdpb_inst_3.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE003F800FFFE1FFF003FFFFFC003FF00F01FE;
defparam sdpb_inst_3.INIT_RAM_25 = 256'hFFFFFFFFFFFFFC001FFFF800000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_26 = 256'h0FFE01FFF83FFE01FFFFFF000FFF03C01FFFE000F8F00707FFFFFFFFFFFFC01F;
defparam sdpb_inst_3.INIT_RAM_27 = 256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam sdpb_inst_3.INIT_RAM_28 = 256'h7001FFF0001FF801C7FFFFFFFFFFFFE003FFFFFFFFFFFFFFC007FFFF00000000;
defparam sdpb_inst_3.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE003FFE03FFE07FF83FFFFFFE001E7F0;
defparam sdpb_inst_3.INIT_RAM_2A = 256'hF800FFFFFFFFFFFFFFF001FFFFE0000000000000003FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2B = 256'hFFF000FFF803FF80FFC1FFFFFFFE007C7F1E001FF00007FC007BFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2D = 256'h0F0FE78003F80001FC001FFFFFFFFFFFFFFE003FFFFFFFFFFFFFFC007FFFFC00;
defparam sdpb_inst_3.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FF003FE00FD07FFFFFFFC0;
defparam sdpb_inst_3.INIT_RAM_2F = 256'hFFFFFF801FFFFFFFFFFFFFFF800FFFFF80000000008000003FFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_30 = 256'hFFFFFFFF80007FC003E000001FFFFFFFFC03C0FFE0003E00007E0007FFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_31 = 256'hFFF00000000500000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_32 = 256'hFFFFC0F00FF8000F80001F8001FFFFFFFFFFFFFFE007FFFFFFFFFFFFFFF001FF;
defparam sdpb_inst_3.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003F80000000007FFFF;
defparam sdpb_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFC00FFFFFFFFFFFFFFFC007FFFFE00000004000000007FFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFF80003F0000000003FFFFFFFFFC1E00FF0001F0000FC0007FFF;
defparam sdpb_inst_3.INIT_RAM_36 = 256'h001FFFFFC00000020000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_37 = 256'hFFFFFFFFFFC7800FC0007C0007F0003FFFFFFFFFFFFFFF801FFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000;
defparam sdpb_inst_3.INIT_RAM_39 = 256'h1FFFFFFFFFFFFFFFE007FFFFFFFFFFFFFFC007FFFFF80000000000000000FFFF;
defparam sdpb_inst_3.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFF00000000000003FFFFFFFFFFDE000F8001F0007FC00;
defparam sdpb_inst_3.INIT_RAM_3B = 256'hFFFFF003FFFFFF00000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3C = 256'h00000FFFFFFFFFFFFC001F8007C003EF800FFFFFFFFFFFFFFFF001FFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000;
defparam sdpb_inst_3.INIT_RAM_3E = 256'hE3E00FFFFFFFFFFFFFFFFC007FFFFFFFFFFFFFFC00FFFFFFE000000000000000;
defparam sdpb_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000003FFFFFFFFFFFF0007F801F003;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_19}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b1;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFF003FFFFFFC20000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_01 = 256'h0000000001FFFFFFFFFFFFC000FF803E01F07807FFFFFFFFFFFFFFFF800FFFFF;
defparam sdpb_inst_4.INIT_RAM_02 = 256'h0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_4.INIT_RAM_03 = 256'h0F80F81E03FFFFFFFFFFFFFFFFE001FFFFFFFFFFFFFF800FFFFFFF8000000000;
defparam sdpb_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000007FFFFFFFFFFFF8003DF0;
defparam sdpb_inst_4.INIT_RAM_05 = 256'h3FFFFFFFFFFFFFE003FFFFFFF00000000000000001FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_06 = 256'hFFF8000000000007FFFFFFFFFFFF800F1F03E0FC0781FFFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_4.INIT_RAM_07 = 256'h0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_08 = 256'h03E1F0F87C01E1FFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFF800FFFFFFFC0000;
defparam sdpb_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000006FFFFFFFFFFFFF8;
defparam sdpb_inst_4.INIT_RAM_0A = 256'hFFF001FFFFFFFFFFFFF8003FFFFFFF80000000000000000FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0B = 256'hFFFFFFFFF000000000007FFFFFFFFFFFFF80781F3E3E0078FFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0C = 256'hF00000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0D = 256'hFFFFF81E03F7FF001E7FFFFFFFFFFFFFFFFFFC007FFFFFFFFFFFF8001FFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0F = 256'hFFFFFFFF001FFFFFFFFFFFFE000FFFFFFFFE00000000000000003FFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFF7F800000000FFFFFFFFFFFFFF07C03FFF8007FFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_11 = 256'hFFFFFF00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFF0F003FF8000FFFFFFFFFFFFFFFFFFFFE001FFFFFFFFFFFF0007FF;
defparam sdpb_inst_4.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000001FFF;
defparam sdpb_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFF8001FFFFFFFFFFFC003FFFFFFFFC00000000000000003FFFFFF;
defparam sdpb_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFE0000000003FFFFFFFFFFFFFF3C003FC0003FFFFFFF;
defparam sdpb_inst_4.INIT_RAM_16 = 256'h00FFFFFFFFF000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_17 = 256'h007FFFFFFFFFFFFFFF0003F0000FFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFE0;
defparam sdpb_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
defparam sdpb_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFE0007FFFFFFFF800000000000000001F;
defparam sdpb_inst_4.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000001FFFFFFFFFFFFFFFE0007C0007FF;
defparam sdpb_inst_4.INIT_RAM_1B = 256'hFFF0003FFFFFFFFE000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1C = 256'h00000003FFFFFFFFFFFFFFF8001F0003FFFFFFFFFFFFFFFFFFFFFC003FFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1D = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam sdpb_inst_4.INIT_RAM_1E = 256'h03FFFFFFFFFFFFFFFFFFFFFF001FFFFFFFFFF8001FFFFFFFFF80000000000000;
defparam sdpb_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000007FFFFFFFFFFFFFFF0003C0;
defparam sdpb_inst_4.INIT_RAM_20 = 256'hFFFFFF80001FFFFFFFFFE000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_21 = 256'hFE00000000001FFFFFFFFFFFFFFFE000F001FFFFFFFFFFFFFFFFFFFFFFE003FF;
defparam sdpb_inst_4.INIT_RAM_22 = 256'h000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_23 = 256'h003C00FFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFC0000FFFFFFFFFF800000000;
defparam sdpb_inst_4.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000003FFFFFFFFFFFFFFFE;
defparam sdpb_inst_4.INIT_RAM_25 = 256'h0007FFFFFFE00003FFFFFFFFFF000000000000000003FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_26 = 256'hFFFFFFC000000000007FFFFFFFFFFFFFFFE00F807FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_27 = 256'h00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_28 = 256'hFFFFFE03E07FFFFFFFFFFFFFFFFFFFFFFFE000FFFFFF300001FFFFFFFFFFC000;
defparam sdpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000001FFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2A = 256'hFFFFFC003FFFFF000000FFFFFFFFFFF800000000000000003FFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2B = 256'hFFFFFFFFFFFC000000000007FFFFFFFFFFFFFFFFE0783FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2C = 256'hFE00000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFC1E1FFFFFFFFFFFFFFFFFFFFFFFFF000C3FFF800000FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000001FFFFFF;
defparam sdpb_inst_4.INIT_RAM_2F = 256'hFFFFFFFFFFC00003C0400007FFFFFFFFFFFFC00000000000000007FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFC000000000003FFFFFFFFFFFFFFFFFC78FFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_31 = 256'hFFFFFFF00000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFF8000060000003FFFFFF;
defparam sdpb_inst_4.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000001F;
defparam sdpb_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFE000000000001FFFFFFFFFFFFFE00000000000000007FFFFF;
defparam sdpb_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFFFFC0000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_37 = 256'h0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000003FF;
defparam sdpb_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000;
defparam sdpb_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFC000000200FFFFFFFFFFFFFFFF8000020000000000F;
defparam sdpb_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000001FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3B = 256'h07FFFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3C = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000C;
defparam sdpb_inst_4.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_4.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000383FFFFFFFFFFFFFFFFE00000000000;
defparam sdpb_inst_4.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_20}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b1;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFF8000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_01 = 256'hFFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam sdpb_inst_5.INIT_RAM_02 = 256'h000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0782FFFFFFFFFFFFFFFFFFFF800000;
defparam sdpb_inst_5.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_06 = 256'hFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_07 = 256'h00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_5.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000003FFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0B = 256'hFFFFFFFFFFFFF80000001E3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0C = 256'hFFFFF80000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000003F8FFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000001FFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFE0001FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_11 = 256'hFFFFFFFFFFF00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF03FFFFF7F;
defparam sdpb_inst_5.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000FFFFF;
defparam sdpb_inst_5.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFF0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_17 = 256'hFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_18 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF;
defparam sdpb_inst_5.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000;
defparam sdpb_inst_5.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FF807FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1C = 256'hFFFFF003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1D = 256'h000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0400;
defparam sdpb_inst_5.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3001FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_21 = 256'hFFFFFFFF0200FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_22 = 256'hFC5000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE061FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_26 = 256'hFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_27 = 256'hFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01EFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000007FFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2C = 256'hFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000002FFFFFFF;
defparam sdpb_inst_5.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFF8100000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3F;
defparam sdpb_inst_5.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007FFFFFFFFFFFFFFFFFFF8200000003F;
defparam sdpb_inst_5.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_36 = 256'h0181FFFFFFFFFFFFFFFFFFFF020000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_5.INIT_RAM_38 = 256'h4000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFE00000;
defparam sdpb_inst_5.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3B = 256'hFFFF00007FFFFFFFFFFFFFFFFFFFFC10000000BFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3D = 256'h8300000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC003FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_21}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b1;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'hFFFFFFF9383FFFFFFFFFFFFFFFFFFFFFFFF0604000007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_02 = 256'hFFFFFE1C8000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE4FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_05 = 256'hFFFFFFFFFF13FFFFFFFFFFFFFFFFFFFFFFFFFFFFC100010001FFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFF0C00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_07 = 256'hFFFFFFFFFFF8600000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF90FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7001FFF;
defparam sdpb_inst_6.INIT_RAM_0A = 256'hFFFFFFFFFFFF10FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0A0200000FFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF38381FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFE080000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0D = 256'hE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF087FFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDE1;
defparam sdpb_inst_6.INIT_RAM_0F = 256'hFFFFFFFFFFFFFE007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC100002001FFF;
defparam sdpb_inst_6.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF870701FFFFFFFFFFFFF0003FFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFF8400000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_12 = 256'hFE3C3C0FFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_13 = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_14 = 256'hFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0800000;
defparam sdpb_inst_6.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1E1E03FFFFFFFFFFFF0000003FFF;
defparam sdpb_inst_6.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_17 = 256'hFFFFFFCF0F007FFFFFFFFFFF80000003FFFFFFFFFFFFFFF807FFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_18 = 256'h00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_19 = 256'h001FFFFFFFFFFFFFE03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sdpb_inst_6.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3C7803FFFFFFFFFFFC00000;
defparam sdpb_inst_6.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8400000003FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1C = 256'hFFFFFFFFFFE1E3C03FFFFFFFFFFFE000000003FFFFFFFFFFFF81FFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1D = 256'hFFFE0C0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1E = 256'h000000007FFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F1F01FFFFFFFFFFFF8;
defparam sdpb_inst_6.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFE387807FFFFFFFFFFFC000000000FFFFFFFFFFC1FFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_22 = 256'hFFFFFFFFF8200000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_23 = 256'hFFFF0000000003FFFFFFFFF93FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9E3C01FFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC01FFFFFFFFFFFFFFF0400000003FFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFE31E20FFFFFFFFFFFFC000000000FFFFFFFFF3FFFFFF;
defparam sdpb_inst_6.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFE000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_28 = 256'hFFFFFFFFF0000000003FFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00007;
defparam sdpb_inst_6.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00F00FFFF;
defparam sdpb_inst_6.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFC0000007F800000001FFFFFFFFFFFFFFFC180800001FFFFF;
defparam sdpb_inst_6.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC01007FFFFFFFFFFFFC000000000FFFFFFFC3FF;
defparam sdpb_inst_6.INIT_RAM_2C = 256'h000FFFFFFFFFFFFFFFFF8200000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2D = 256'h0FFFFFFFFFFFFF0000000003FFFFFF87FFFFFFFFFFFFFFFFF000000000000000;
defparam sdpb_inst_6.INIT_RAM_2E = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000;
defparam sdpb_inst_6.INIT_RAM_2F = 256'h8FFFFFFFFFFFFFFFFC000FFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFF080000000;
defparam sdpb_inst_6.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFC000000000FFFFFF;
defparam sdpb_inst_6.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0800000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_32 = 256'hC70003FFFFFFFFFFFFF0000000007FFFFF0FFFFFFFFFFFFFFFC003FFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_33 = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_34 = 256'hFFFF1FFFFFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC200;
defparam sdpb_inst_6.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03807FFFFFFFFFFFFFE000000003F;
defparam sdpb_inst_6.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8400000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_37 = 256'hFFFFF00103FFFFFFFFFFFFFF800000000FFFFF1FFFFFFFFFFFFFF807FFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_38 = 256'hFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_39 = 256'h0007FFFE3FFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFE00000;
defparam sdpb_inst_6.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3C = 256'hFFFFFFFFFE0001FFFFFFFFFFFFFFFC00000003FFFE3FFFFFFFFFFFFFE07FFFFF;
defparam sdpb_inst_6.INIT_RAM_3D = 256'hFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3E = 256'h00000001FFFE3FFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFF;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_22}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b1;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFE0000001FFFE3FFFFFFFFFFFFFC1FF;
defparam sdpb_inst_7.INIT_RAM_02 = 256'hFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_03 = 256'hFFFFF8000000FFFE3FFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_05 = 256'h83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFF;
defparam sdpb_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFF0000007FFF3FFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_08 = 256'hFFFFFFFFFFC000003FFF3FFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFF;
defparam sdpb_inst_7.INIT_RAM_0A = 256'hFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001F;
defparam sdpb_inst_7.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFF800003FFF1FFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFE00001FFF1FFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0E = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FF;
defparam sdpb_inst_7.INIT_RAM_0F = 256'hFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000;
defparam sdpb_inst_7.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFC0001FFF8FFFFF;
defparam sdpb_inst_7.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_12 = 256'h003FFFFFFFFFFFFFFFFFF8001FFF8FFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_13 = 256'h8000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sdpb_inst_7.INIT_RAM_14 = 256'hFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFF001FFFCF;
defparam sdpb_inst_7.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_17 = 256'hFFF0000FFFFFFFFFFFFFFFFFFFC01FFFC7FFFFFFFFFFFC1FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_18 = 256'hFFFFFE0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_19 = 256'hFFE7FFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFC3F;
defparam sdpb_inst_7.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1C = 256'hFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFF83FFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1D = 256'hFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1E = 256'hFFFFFFF9FFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000100001FFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_21 = 256'hFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFF87FFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFE0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_23 = 256'hFFFFFFFFFFFEFFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FF;
defparam sdpb_inst_7.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFF87FFFFF;
defparam sdpb_inst_7.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFBFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_29 = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam sdpb_inst_7.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFF87F;
defparam sdpb_inst_7.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000200003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2E = 256'h000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFF;
defparam sdpb_inst_7.INIT_RAM_2F = 256'hFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sdpb_inst_7.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_32 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_33 = 256'hFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam sdpb_inst_7.INIT_RAM_34 = 256'hFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFEFFFF;
defparam sdpb_inst_7.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003FFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_37 = 256'hE00007FFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_38 = 256'hFFFFFFFFFC0000400007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_39 = 256'h9FFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3C = 256'hFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF8FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3E = 256'hFFFFE7FFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[30:0],sdpb_inst_8_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_23}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_8.READ_MODE = 1'b1;
defparam sdpb_inst_8.BIT_WIDTH_0 = 1;
defparam sdpb_inst_8.BIT_WIDTH_1 = 1;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_8.RESET_MODE = "SYNC";
defparam sdpb_inst_8.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003FFFF;
defparam sdpb_inst_8.INIT_RAM_01 = 256'hFFFFFFFFFF00003FFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFE3FFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFC0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_03 = 256'hFFFFFFFFFDFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_04 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001FFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000;
defparam sdpb_inst_8.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF8FFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_08 = 256'hFFFFFFFFFFFFFF3FFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_09 = 256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003FFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam sdpb_inst_8.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFE3FFFFF;
defparam sdpb_inst_8.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFE7FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0E = 256'hFF80000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFF;
defparam sdpb_inst_8.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFCF;
defparam sdpb_inst_8.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000080000FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_13 = 256'hFFFFFFFE0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001F;
defparam sdpb_inst_8.INIT_RAM_14 = 256'hFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFFFFFCFFFFFF;
defparam sdpb_inst_8.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000003FFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_17 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_18 = 256'hFFFFFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sdpb_inst_8.INIT_RAM_19 = 256'hFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFF9F;
defparam sdpb_inst_8.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000FFFFFF;
defparam sdpb_inst_8.INIT_RAM_1C = 256'hFFF80000FFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFE0000100001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1E = 256'hFFE7FFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000003;
defparam sdpb_inst_8.INIT_RAM_21 = 256'hFFFFFFFE00001FFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFC7FFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_23 = 256'hFFFFFFFDFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_24 = 256'h000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000;
defparam sdpb_inst_8.INIT_RAM_26 = 256'hFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF9FFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_28 = 256'hFFFFFFFFFFFFBFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_29 = 256'hC0000200001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFE3FFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000003FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFE7FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2E = 256'hFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFC00001FFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFCFFF;
defparam sdpb_inst_8.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_33 = 256'hFFFFFFFFFFFC0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFF;
defparam sdpb_inst_8.INIT_RAM_34 = 256'hF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC000007FFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFF;
defparam sdpb_inst_8.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000003FFFFFFF;
defparam sdpb_inst_8.INIT_RAM_37 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000;
defparam sdpb_inst_8.INIT_RAM_39 = 256'hFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFCFFF;
defparam sdpb_inst_8.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FF;
defparam sdpb_inst_8.INIT_RAM_3C = 256'h8000007FFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFC0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3E = 256'hF9FFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3F = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000001FFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[30:0],sdpb_inst_9_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_24}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_9.READ_MODE = 1'b1;
defparam sdpb_inst_9.BIT_WIDTH_0 = 1;
defparam sdpb_inst_9.BIT_WIDTH_1 = 1;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_9.RESET_MODE = "SYNC";
defparam sdpb_inst_9.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000;
defparam sdpb_inst_9.INIT_RAM_01 = 256'hFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFE3FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_03 = 256'hFFFFFF7FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_04 = 256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sdpb_inst_9.INIT_RAM_06 = 256'hFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFCFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_08 = 256'hFFFFFFFFFFE7FFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_09 = 256'hFFFF80000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_0B = 256'hFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFF9FFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000003FFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFCFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_0E = 256'hFFFFFFFFFE00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFC000003FFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFF3FFFF;
defparam sdpb_inst_9.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000FFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFF9FFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFF80000000001FFFFFFFFFFFFFFFFFFFFFFFFFE000000FFFFF7;
defparam sdpb_inst_9.INIT_RAM_14 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFE0000007FFFFCFFFFFFFFFFFFFFFFFFFFE7FFFFFFFE;
defparam sdpb_inst_9.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000003FFF;
defparam sdpb_inst_9.INIT_RAM_17 = 256'hFFFF1FFFFFFFFFFFFFFFFFFFF3FFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFE00000000007FFFFFFFFFFFFFFFFFFFFFFFF0000003F;
defparam sdpb_inst_9.INIT_RAM_19 = 256'hFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_1A = 256'h00FFFFFFFFFFFFFFFFFFFFFFFF0000000FFFFFE7FFFFFFFFFFFFFFFFFFFCFFFF;
defparam sdpb_inst_9.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000;
defparam sdpb_inst_9.INIT_RAM_1C = 256'h0001FFFFF8FFFFFFFFFFFFFFFFFFFE7FFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF80000000001FFFFFFFFFFFFFFFFFFFFFFF8000;
defparam sdpb_inst_9.INIT_RAM_1E = 256'h9FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_1F = 256'h00000003FFFFFFFFFFFFFFFFFFFFFFC00000007FFFFE3FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_20 = 256'hFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam sdpb_inst_9.INIT_RAM_21 = 256'hF00000000FFFFF87FFFFFFFFFFFFFFFFFFE7FFFFFFFC7FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000007FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_23 = 256'hFFFFF3FFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_24 = 256'hFFC0000000000FFFFFFFFFFFFFFFFFFFFFF800000003FFFFE1FFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_26 = 256'hFFFFFE00000000FFFFF87FFFFFFFFFFFFFFFFFFCFFFFFFFF8FFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000001FFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_28 = 256'hFFFFFFFFFE7FFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_29 = 256'hFFFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFF800000003FFFFE1FFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2B = 256'hFFFFFFFFFFC00000000FFFFF87FFFFFFFFFFFFFFFFFF9FFFFFFFF9FFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFE7FFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FFFFFF;
defparam sdpb_inst_9.INIT_RAM_2E = 256'hFFFFFFFFFFFFFC0000100003FFFFFFFFFFFFFFFFFE0FF000000007FFFFC3FFFF;
defparam sdpb_inst_9.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_30 = 256'hFFFFFFFFFFFF03FC00000001FFFFF0FFFFFFFFFFFFFFFFFFF1FFFFFFFF3FFFFF;
defparam sdpb_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFF;
defparam sdpb_inst_9.INIT_RAM_32 = 256'h3FFFFFFFFFFFFFFFFFFCFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07F;
defparam sdpb_inst_9.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFE87F00000000FFFFF8;
defparam sdpb_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFF1FE00000003FFFFC0FFFFFFFFFFFFFFFFFFF3FFFFFFFE3;
defparam sdpb_inst_9.INIT_RAM_36 = 256'hF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000F;
defparam sdpb_inst_9.INIT_RAM_37 = 256'hFFFF07FFFFFFFFFFFFFFFFFFDFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFF4FF80000001F;
defparam sdpb_inst_9.INIT_RAM_39 = 256'hFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFFFFFFFFFF0000000FFFFF83FFFFFFFFFFFFFFFFFFE7FFFF;
defparam sdpb_inst_9.INIT_RAM_3B = 256'hFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000;
defparam sdpb_inst_9.INIT_RAM_3C = 256'h0007FFFFC0FFFFFFFFFFFFFFFFFFF9FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000003FFFFFFFFFFFFFFFFFFFFFC000;
defparam sdpb_inst_9.INIT_RAM_3E = 256'h7FFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3F = 256'hE00000000FFFFFFFFFFFFFFFFFFFFFF8000003FFFFE07FFFFFFFFFFFFFFFFFFE;

SDPB sdpb_inst_10 (
    .DO({sdpb_inst_10_dout_w[30:0],sdpb_inst_10_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_25}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_10.READ_MODE = 1'b1;
defparam sdpb_inst_10.BIT_WIDTH_0 = 1;
defparam sdpb_inst_10.BIT_WIDTH_1 = 1;
defparam sdpb_inst_10.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_10.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_10.RESET_MODE = "SYNC";
defparam sdpb_inst_10.INIT_RAM_00 = 256'hFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_01 = 256'hFF800003FFFFF03FFFFFFFFFFFFFFFFFFF9FFFFFFFF1FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000007FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_03 = 256'hFFFFCFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_04 = 256'hFFFFFFC0000001FFFFFFFFFFFFFFFFF7FFFFF00003FFFFE00FFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_06 = 256'hF9FFFFFF8003FFFFF807FFFFFFFFFFFFFFFFFFF3FFFFFFFF3FFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_08 = 256'hFFFFFFFFFCFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_09 = 256'hFFFFFFFFFFFF8000007FFFFFFFFFFFFFFFF97FFFFFFF7FFFFFF803FFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0B = 256'hFFFFFE7FFFFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFF3FFFFFFFF3FFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800003FFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFCFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFBFF;
defparam sdpb_inst_10.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFF88003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00FFFFFF;
defparam sdpb_inst_10.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFC3FFFFFFDFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE007FFFFFFFFFFFFFFFFFFFE7FFFFFFFF3FFFFF;
defparam sdpb_inst_10.INIT_RAM_11 = 256'hFF03FFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07FFFFFFF;
defparam sdpb_inst_10.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFF9FFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF;
defparam sdpb_inst_10.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFFFF003F;
defparam sdpb_inst_10.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFF803FFFFFE3FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFE00FFFFFFFFFFFFF001FFFFFFFFFFFFFFFFFFFFE7FFFFFFFE3;
defparam sdpb_inst_10.INIT_RAM_16 = 256'hFFFFFFC003FFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_17 = 256'h801FFFFFFFFFFFFFFFFFFFFF3FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFE7;
defparam sdpb_inst_10.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE003FFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_19 = 256'hFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFE0007FFFFF03FFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFFE00FFFFFFFFFFFFFFFFFFFFFCFFFFF;
defparam sdpb_inst_10.INIT_RAM_1B = 256'hFFFCFFFFFFF00007FFFFC03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1C = 256'hFFFFF807FFFFFFFFFFFFFFFFFFFFF7FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFCF;
defparam sdpb_inst_10.INIT_RAM_1E = 256'hFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFC00007FFFF007FFFFFF;
defparam sdpb_inst_10.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFE7FFFFFC03FFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_10.INIT_RAM_20 = 256'hFFFFFFFF3FFFFFFE000007FFFE007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_21 = 256'hFFF3FFFFFF01FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF9FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0083FF;
defparam sdpb_inst_10.INIT_RAM_23 = 256'hFFFF9FFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFD8FFFFFFF0000007FFF8007;
defparam sdpb_inst_10.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFA00001FFFFC7FFDFFC0FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_25 = 256'hFFFFFFFFFFFFE7FFFFFF80000007FFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_26 = 256'h000FFFFF0FFE7FE07FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF3FFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_27 = 256'hFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400;
defparam sdpb_inst_10.INIT_RAM_28 = 256'hFFFFFFFFFBFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFB1FFFFFFC0000000FF;
defparam sdpb_inst_10.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFF000000FFFFC1FFBFF81FFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFDCFFFFFFF00000000FFFC0003FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2B = 256'hFF0000001FFFF80FC7FE0FFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFF3FFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2C = 256'h0000FFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F;
defparam sdpb_inst_10.INIT_RAM_2D = 256'hFFFFFFFFFFFFFF3FFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFF80000;
defparam sdpb_inst_10.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFF80000003FFF80079FF83FFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFB9FFFFFFC000000000FFFC0001FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_30 = 256'hFFE1FFC00000041FF800003FF0FFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFE7FFFFF;
defparam sdpb_inst_10.INIT_RAM_31 = 256'h0000000000FFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFF7FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFF;
defparam sdpb_inst_10.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF03FC01C000061FE000007FC3FFF;
defparam sdpb_inst_10.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF607FFFFF80000000000FFFC0001FFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_35 = 256'hFFFFFFFC07C00F0000020F800003FF0FFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFE7;
defparam sdpb_inst_10.INIT_RAM_36 = 256'hFFFFC00000000000FFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_37 = 256'h83FFFFFFFFFFFFFFFFFFFFFF7FFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFF81F;
defparam sdpb_inst_10.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00400FC0000030400000FF;
defparam sdpb_inst_10.INIT_RAM_39 = 256'hFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFEC07FFFFE000000000000FFFC000FFFFFF;
defparam sdpb_inst_10.INIT_RAM_3A = 256'hFFFFFFFFFFFF80000FF00000018000003FE0FFFFFFFFFFFFFFFFFFFFFF9FFFFF;
defparam sdpb_inst_10.INIT_RAM_3B = 256'hFE03FFFFF8000000000001FFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3C = 256'h001FF83FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00007FC0000000800;
defparam sdpb_inst_10.INIT_RAM_3E = 256'hFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFD80FFFFFC0000000000003FFFC001;
defparam sdpb_inst_10.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFF00003FE00000000000003FF0FFFFFFFFFFFFFFFFFFFFFF9;

SDPB sdpb_inst_11 (
    .DO({sdpb_inst_11_dout_w[30:0],sdpb_inst_11_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_26}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_11.READ_MODE = 1'b1;
defparam sdpb_inst_11.BIT_WIDTH_0 = 1;
defparam sdpb_inst_11.BIT_WIDTH_1 = 1;
defparam sdpb_inst_11.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_11.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_11.RESET_MODE = "SYNC";
defparam sdpb_inst_11.INIT_RAM_00 = 256'hFFFFFF607FFFFE0000000000001FFFFA001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_01 = 256'h00000000FF83FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFE3FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_02 = 256'hFF8141FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FF800000;
defparam sdpb_inst_11.INIT_RAM_03 = 256'hFFFF9FFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFB01FFFFF0000000000000FFF;
defparam sdpb_inst_11.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFF00007FC00000000000001FE0FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_05 = 256'hFFFFFFFFFFEC0FFFFFC0000000000003FFFFF85C1FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_06 = 256'h00000000000007F83FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFE7FFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_07 = 256'h01FFFFFF89C1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007F0;
defparam sdpb_inst_11.INIT_RAM_08 = 256'hFFFFFFFFFBFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFF603FFFFE00000000000;
defparam sdpb_inst_11.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE000007800000000000001FC0FFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFD81FFFFFF000000000000FFFFFFFC783FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0B = 256'h0004000000418000003F83FFFFFFFFFFFFFFFFFFFFFCFFFFFFFFC7FFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0C = 256'h0000003FFFFFFF8383FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800;
defparam sdpb_inst_11.INIT_RAM_0D = 256'hFFFFFFFFFFFFFF3FFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFF607FFFFFF00000;
defparam sdpb_inst_11.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000001FF8000007C0FFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFD03FFFFFFF80000000001FFFFFFFF8303FFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_10 = 256'hFF80000000000003FC000000F03FFFFFFFFFFFFFFFFFFFFFCFFFFFFFFCFFFFFF;
defparam sdpb_inst_11.INIT_RAM_11 = 256'hF8000000000FFFFFFFFF8303FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFF3FFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFF41FFFFFFF;
defparam sdpb_inst_11.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000007F0000001C0FFF;
defparam sdpb_inst_11.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFD07FFFFFFFF8000000003FFFFFFFFF8103FFFFF;
defparam sdpb_inst_11.INIT_RAM_15 = 256'hFFFFFFFC000000000000078000000207FFFFFFFFFFFFFFFFFFFFFCFFFFFFFF9F;
defparam sdpb_inst_11.INIT_RAM_16 = 256'hFFFFFFFC00000001FFFFFFFFFFC103FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_17 = 256'h01FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFBFF;
defparam sdpb_inst_11.INIT_RAM_18 = 256'h3FF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000040000000;
defparam sdpb_inst_11.INIT_RAM_19 = 256'hFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000FFFFFFFFFFFC00;
defparam sdpb_inst_11.INIT_RAM_1A = 256'hFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFF9FFFFF;
defparam sdpb_inst_11.INIT_RAM_1B = 256'hFFFFFFFFFFFFFC0000003FFFFFFFFFFFC007FC3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1C = 256'h0000001FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1D = 256'hFFFE007F0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000;
defparam sdpb_inst_11.INIT_RAM_1E = 256'hFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000001FFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFE00000000000000000000000FFFFFFFFFFFFFFFFFFFFFF9;
defparam sdpb_inst_11.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFF00403FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_21 = 256'h000000000003FFFFFFFFFFFFFFFFFFFFFCFFFFFFFF8FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_22 = 256'hFFFFFFFFEF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000;
defparam sdpb_inst_11.INIT_RAM_23 = 256'hFFFF3FFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFF;
defparam sdpb_inst_11.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFF87C003FFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_26 = 256'h00000000000000007FFFFFFFFFFFFFFFFFFFFFCFFFFFFFF9FFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_27 = 256'hFFFFFFFFFFFFFE03E00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000;
defparam sdpb_inst_11.INIT_RAM_28 = 256'hFFFFFFFFF3FFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam sdpb_inst_11.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000001FFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE007FFFFFFFFFFFFF001E01FFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2B = 256'h000000000000000003800FFFFFFFFFFFFFFFFFFFFFF9FFFFFFFF3FFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2C = 256'hFFF01FFFFFFFFFFFFFC001F01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam sdpb_inst_11.INIT_RAM_2D = 256'hFFFFFFFFFFFFFE7FFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000007003FFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFF0000F83FFFF;
defparam sdpb_inst_11.INIT_RAM_30 = 256'hFFFF8000000000000000001E01FFFFFFFFFFFFFFFFFFFFFF9FFFFFFFE3FFFFFF;
defparam sdpb_inst_11.INIT_RAM_31 = 256'hFFFFFFFFFBFFFFFFFFFFFFF800007C7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFE7FFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000C2007FFF;
defparam sdpb_inst_11.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000003;
defparam sdpb_inst_11.INIT_RAM_35 = 256'hFFFFFFFFFF000000000000000038003FFFFFFFFFFFFFFFFFFFFFF3FFFFFFFC7F;
defparam sdpb_inst_11.INIT_RAM_36 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFF8000001F7FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_37 = 256'h1FFFFFFFFFFFFFFFFFFFFFFDFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam sdpb_inst_11.INIT_RAM_38 = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000800000000000700;
defparam sdpb_inst_11.INIT_RAM_39 = 256'hFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sdpb_inst_11.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFE000180000000003C0007FFFFFFFFFFFFFFFFFFFFFF3FFFFF;
defparam sdpb_inst_11.INIT_RAM_3B = 256'hFFFF047FFFFFFFFFDFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3C = 256'h6D0003FFFFFFFFFFFFFFFFFFFFFF8FFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3D = 256'hFFF800000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000CE30000000;
defparam sdpb_inst_11.INIT_RAM_3E = 256'hFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007FFFFFFFF01FFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFE0017DDC000007B0001FFFFFFFFFFFFFFFFFFFFFFE7;

SDPB sdpb_inst_12 (
    .DO({sdpb_inst_12_dout_w[30:0],sdpb_inst_12_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_27}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_12.READ_MODE = 1'b1;
defparam sdpb_inst_12.BIT_WIDTH_0 = 1;
defparam sdpb_inst_12.BIT_WIDTH_1 = 1;
defparam sdpb_inst_12.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_12.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_12.RESET_MODE = "SYNC";
defparam sdpb_inst_12.INIT_RAM_00 = 256'hFFFFFFFFFC007FFFFFFC001FFFFFFFFFFFFFFE000000007FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_01 = 256'h1819C60000FFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFE7FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_02 = 256'hFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001EFC0;
defparam sdpb_inst_12.INIT_RAM_03 = 256'hFFF87FFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00FFFFFF80001FFFFFF;
defparam sdpb_inst_12.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC000360E686F000007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFF084FFFFE000001FFFFFFFFFFFFFC000000003FFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_06 = 256'h00002DF18C00007FFFFFFFFFFFFFFFFFFFFFFC07FFFFFFCFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_07 = 256'hFFFFFFFFFFFFE000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sdpb_inst_12.INIT_RAM_08 = 256'hFFFFFFFF01FFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE287FFFF8000001;
defparam sdpb_inst_12.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000003786000003FFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFC1E1FFFF8000001FFFFFFFFFFFF8000000003FFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0B = 256'hFFFFE00000000000001FFFFFFFFFFFFFFFFFFFFFFFC07FFFFFF8FFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0C = 256'h000001FFFFFFFFFFFC0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0D = 256'hFFFFFFFFFFFFE03FFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8443FFFF0;
defparam sdpb_inst_12.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000001FFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF8407FFFF0000001FFFFFFFFFFF0000000001FF;
defparam sdpb_inst_12.INIT_RAM_10 = 256'hFFFFFFFFFFF000000000001FFFFFFFFFFFFFFFFFFFFFFFF80FFFFFFF1FFFFFFF;
defparam sdpb_inst_12.INIT_RAM_11 = 256'h7FFFF0000001BFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFE03FFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA00;
defparam sdpb_inst_12.INIT_RAM_13 = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000001FFFFFFF;
defparam sdpb_inst_12.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0AFFFFE00000007FFFFFFFFC0000000;
defparam sdpb_inst_12.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFFFFFF81FFFFFFE3FF;
defparam sdpb_inst_12.INIT_RAM_16 = 256'hFFF011FFFFE00000007FFFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFC07FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_18 = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01000003FFF;
defparam sdpb_inst_12.INIT_RAM_19 = 256'hFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003FFFFE00000007FFFFFFF800;
defparam sdpb_inst_12.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFF01FFFFF;
defparam sdpb_inst_12.INIT_RAM_1B = 256'hFFFFFFFFF807FFFFE00000007FFFFFFC00000000003FFF9FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1D = 256'hFF00000000000FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC007;
defparam sdpb_inst_12.INIT_RAM_1E = 256'hFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFE00000007FFFF;
defparam sdpb_inst_12.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03;
defparam sdpb_inst_12.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFCFFFFFFC0000000FFFFFF800000000003FFFD3FFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80FFFFFF81FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_22 = 256'h0FFFFFC00000000000FFFE67FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_23 = 256'hFFE07FFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFC000000;
defparam sdpb_inst_12.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFC73FFFFC0000000FFFFE000000000003FFF9CFFFFFF;
defparam sdpb_inst_12.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01FFFFFF81FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_27 = 256'h0000001FFFF000000000000FFFF79FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_28 = 256'hFFFFFFFC07FFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC73FFFFC;
defparam sdpb_inst_12.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFCF3FFFF80000001FFF8000000000003FFFDFF;
defparam sdpb_inst_12.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01FFFFFF03FFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2C = 256'hBFFFF00000003FFC000000000000FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2D = 256'hFFFFFFFFFFFF80FFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F;
defparam sdpb_inst_12.INIT_RAM_2E = 256'hFFDFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1F3FFFF00000007FE0000000000007F;
defparam sdpb_inst_12.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FFFFFF03FFFFFFF;
defparam sdpb_inst_12.INIT_RAM_31 = 256'hFFFE3F3FFFF0000000FF0000000000001FFFF7FDFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFF80FFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_33 = 256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3F3FFFF0000001F8000000000;
defparam sdpb_inst_12.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFF03FF;
defparam sdpb_inst_12.INIT_RAM_36 = 256'hFFFFFFFFFFFF3FFFFC000001C0000000000003FFFF7FEFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_38 = 256'h00000000FFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_39 = 256'hE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFC00000300000;
defparam sdpb_inst_12.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFC0000060000000000007FFFF87FFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3D = 256'hC000000000001FFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3E = 256'hFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFC00000;
defparam sdpb_inst_12.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_13 (
    .DO({sdpb_inst_13_dout_w[30:0],sdpb_inst_13_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_28}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_13.READ_MODE = 1'b1;
defparam sdpb_inst_13.BIT_WIDTH_0 = 1;
defparam sdpb_inst_13.BIT_WIDTH_1 = 1;
defparam sdpb_inst_13.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_13.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_13.RESET_MODE = "SYNC";
defparam sdpb_inst_13.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFEC07FFFFC00001800000000000FFFFFF87FFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_02 = 256'h800003000000000003FFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_03 = 256'hFFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFFF;
defparam sdpb_inst_13.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFEC0FFFFF80000C00000000001FFFFFFFCFFFF;
defparam sdpb_inst_13.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_07 = 256'h0FFFFF80001800000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFF80FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_13.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FFFFF8000300000000003FFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0C = 256'hFFFFFC1FFFFF800060000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFF0000C0000000007FF;
defparam sdpb_inst_13.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_11 = 256'hFFFFFFFFFFFC3FFFFF00018000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_13 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFF00030000000;
defparam sdpb_inst_13.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFC3FFFFF0006000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_18 = 256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFE000C0;
defparam sdpb_inst_13.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFC7FFFFE00100000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1D = 256'hE0020000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF87FFFF;
defparam sdpb_inst_13.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF87FFFFC0040000003FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_22 = 256'h87FFFB0018000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFE0003000000FFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_27 = 256'hFFFFFF8FFFC000600000FFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFC00080000FFFFFFFF8F;
defparam sdpb_inst_13.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2C = 256'hFFFFFFFFFFFF9FFF00010000FFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2E = 256'hFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFF80706001FFFFFF;
defparam sdpb_inst_13.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFF9FEC7F1C03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFF1FFF;
defparam sdpb_inst_13.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFF;
defparam sdpb_inst_13.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3D = 256'hF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_14 (
    .DO({sdpb_inst_14_dout_w[30:0],sdpb_inst_14_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_29}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_14.READ_MODE = 1'b1;
defparam sdpb_inst_14.BIT_WIDTH_0 = 1;
defparam sdpb_inst_14.BIT_WIDTH_1 = 1;
defparam sdpb_inst_14.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_14.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_14.RESET_MODE = "SYNC";
defparam sdpb_inst_14.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC107FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_02 = 256'hFFFFFFC207FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC801FFFFFFFFCFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_07 = 256'hFFFFFFFFFFFFC001FFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80C1FFFFFFE7FFFFF;
defparam sdpb_inst_14.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFF8181FFFFFE1F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF84E3FFFFF0F;
defparam sdpb_inst_14.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFA48FFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_13 = 256'hFF2FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD005F;
defparam sdpb_inst_14.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800BFFC7FFEFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_18 = 256'hF8013FF8FFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA47FF87FF3FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1D = 256'hFFFFFFFCC0FFF87FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01FFF87F9FFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_22 = 256'hFFFFFFFFFFFFFF07FFFC7DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFF81FFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3F = 256'h000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[17]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clkb),
  .CE(oce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[16]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clkb),
  .CE(oce)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[15]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_5 (
  .Q(dff_q_5),
  .D(dff_q_4),
  .CLK(clkb),
  .CE(oce)
);
DFFE dff_inst_6 (
  .Q(dff_q_6),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_7 (
  .Q(dff_q_7),
  .D(dff_q_6),
  .CLK(clkb),
  .CE(oce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sdpb_inst_2_dout[0]),
  .I1(sdpb_inst_3_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sdpb_inst_4_dout[0]),
  .I1(sdpb_inst_5_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sdpb_inst_6_dout[0]),
  .I1(sdpb_inst_7_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(sdpb_inst_8_dout[0]),
  .I1(sdpb_inst_9_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(sdpb_inst_10_dout[0]),
  .I1(sdpb_inst_11_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sdpb_inst_12_dout[0]),
  .I1(sdpb_inst_13_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_5)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_5)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_5)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_6),
  .I1(sdpb_inst_14_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_3)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_3)
);
MUX2 mux_inst_14 (
  .O(dout[0]),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_1)
);
endmodule //Gowin_SDPB
