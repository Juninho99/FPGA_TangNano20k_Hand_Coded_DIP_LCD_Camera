//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Thu Aug 31 18:45:34 2023

module Gowin_pROM4 (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [16:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [1:1] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [1:1] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [1:1] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [1:1] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [2:2] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [2:2] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [2:2] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [2:2] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [3:3] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [3:3] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [3:3] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [3:3] prom_inst_15_dout;
wire [30:0] prom_inst_16_dout_w;
wire [0:0] prom_inst_16_dout;
wire [30:0] prom_inst_17_dout_w;
wire [1:1] prom_inst_17_dout;
wire [30:0] prom_inst_18_dout_w;
wire [2:2] prom_inst_18_dout;
wire [30:0] prom_inst_19_dout_w;
wire [3:3] prom_inst_19_dout;
wire [29:0] prom_inst_20_dout_w;
wire [1:0] prom_inst_20_dout;
wire [29:0] prom_inst_21_dout_w;
wire [3:2] prom_inst_21_dout;
wire [27:0] prom_inst_22_dout_w;
wire [3:0] prom_inst_22_dout;
wire [30:0] prom_inst_23_dout_w;
wire [4:4] prom_inst_23_dout;
wire [30:0] prom_inst_24_dout_w;
wire [4:4] prom_inst_24_dout;
wire [30:0] prom_inst_25_dout_w;
wire [4:4] prom_inst_25_dout;
wire [30:0] prom_inst_26_dout_w;
wire [4:4] prom_inst_26_dout;
wire [30:0] prom_inst_27_dout_w;
wire [5:5] prom_inst_27_dout;
wire [30:0] prom_inst_28_dout_w;
wire [5:5] prom_inst_28_dout;
wire [30:0] prom_inst_29_dout_w;
wire [5:5] prom_inst_29_dout;
wire [30:0] prom_inst_30_dout_w;
wire [5:5] prom_inst_30_dout;
wire [30:0] prom_inst_31_dout_w;
wire [6:6] prom_inst_31_dout;
wire [30:0] prom_inst_32_dout_w;
wire [6:6] prom_inst_32_dout;
wire [30:0] prom_inst_33_dout_w;
wire [6:6] prom_inst_33_dout;
wire [30:0] prom_inst_34_dout_w;
wire [6:6] prom_inst_34_dout;
wire [30:0] prom_inst_35_dout_w;
wire [7:7] prom_inst_35_dout;
wire [30:0] prom_inst_36_dout_w;
wire [7:7] prom_inst_36_dout;
wire [30:0] prom_inst_37_dout_w;
wire [7:7] prom_inst_37_dout;
wire [30:0] prom_inst_38_dout_w;
wire [7:7] prom_inst_38_dout;
wire [30:0] prom_inst_39_dout_w;
wire [4:4] prom_inst_39_dout;
wire [30:0] prom_inst_40_dout_w;
wire [5:5] prom_inst_40_dout;
wire [30:0] prom_inst_41_dout_w;
wire [6:6] prom_inst_41_dout;
wire [30:0] prom_inst_42_dout_w;
wire [7:7] prom_inst_42_dout;
wire [29:0] prom_inst_43_dout_w;
wire [5:4] prom_inst_43_dout;
wire [29:0] prom_inst_44_dout_w;
wire [7:6] prom_inst_44_dout;
wire [27:0] prom_inst_45_dout_w;
wire [7:4] prom_inst_45_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire dff_q_7;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_0.INIT = 16'h0002;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_1.INIT = 16'h0008;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_2.INIT = 16'h0020;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_3.INIT = 16'h0080;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_4.INIT = 16'h0200;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad[13]),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_5.INIT = 16'h0400;
LUT2 lut_inst_6 (
  .F(lut_f_6),
  .I0(ce),
  .I1(lut_f_5)
);
defparam lut_inst_6.INIT = 4'h8;
LUT5 lut_inst_7 (
  .F(lut_f_7),
  .I0(ad[12]),
  .I1(ad[13]),
  .I2(ad[14]),
  .I3(ad[15]),
  .I4(ad[16])
);
defparam lut_inst_7.INIT = 32'h00400000;
LUT2 lut_inst_8 (
  .F(lut_f_8),
  .I0(ce),
  .I1(lut_f_7)
);
defparam lut_inst_8.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b1;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hBDFAFF8B31EDFD48784B49207C73B37E9FFF0599B371FEB0E060DFFE1403DB3E;
defparam prom_inst_0.INIT_RAM_01 = 256'hBFD97E50D3EF603F7A2FE27A5326F682AE65158005D635B7F0831C68BB02791F;
defparam prom_inst_0.INIT_RAM_02 = 256'h9767EB1BE90F9DEE20EF1BD6069FD7E70B4FDDD0277EE4FF027E811F07CBD7BF;
defparam prom_inst_0.INIT_RAM_03 = 256'h40077B697FF994DAE323F4F7BB7F7FFFDC683FDCC38DE11316E3BFAF42BC6E48;
defparam prom_inst_0.INIT_RAM_04 = 256'hE7CDD3343BDE68780BA6FE41053E0444E22E1490BA99BF89F31787507BC52480;
defparam prom_inst_0.INIT_RAM_05 = 256'h8A45BE84A6F141BD187ED4079ED19C04C07F013839FF98BEB9FFC8197E1D8007;
defparam prom_inst_0.INIT_RAM_06 = 256'h1FC0980EE7FE49AF7F310A3200E001999A74FD14F7AFDE0771C7F9F55101B6AB;
defparam prom_inst_0.INIT_RAM_07 = 256'hE0F870B375B3BB3E01BBBFAA705C9B5AF347C731CC005F4A9EB481E6DE7B0100;
defparam prom_inst_0.INIT_RAM_08 = 256'hFEB6239D23CBA9AE76DFE621E9B0806002021B79DFCE7B4C02CC90896807AB42;
defparam prom_inst_0.INIT_RAM_09 = 256'h2100627DBA1E840007F019E54B66482F42CE07C3BFF6F840BBCEB0571B763F67;
defparam prom_inst_0.INIT_RAM_0A = 256'hBFB000EFFDDE080E4C9656E3E60CF277A4F19B0CDE91B21C79FE13346630204E;
defparam prom_inst_0.INIT_RAM_0B = 256'h8C29C3C3936E429E7F97CAC7F00813F65818FEE807A0C082F8E3DB52D87B88E0;
defparam prom_inst_0.INIT_RAM_0C = 256'h01EF86963030446DFBAC7491CBC0027FB02C0487C78C45DC3453E8CC4E3FE598;
defparam prom_inst_0.INIT_RAM_0D = 256'h34C020ADE378F14AA7DD4E812F99F653E56CC3711774191F0FB09EAA4008B428;
defparam prom_inst_0.INIT_RAM_0E = 256'hDBF9CCB6CA7646414C6713E030EF080063E020880CDD1FCD823B427B800093EE;
defparam prom_inst_0.INIT_RAM_0F = 256'h5E02800150BEF7C1FFE719DE0C3FFFC1A4016B1EFF9D0B450B516644315D8A63;
defparam prom_inst_0.INIT_RAM_10 = 256'h00E2DF656A6C3C7DC3AF2B120001DEE299703A3769984E9DF6B1362C3B00241E;
defparam prom_inst_0.INIT_RAM_11 = 256'hFECDFD03E06647866F8FF7E0140739C786440D0443F3FFAFE2538AEF05FCE8D5;
defparam prom_inst_0.INIT_RAM_12 = 256'h910F8110FEFFE5F94162ADC17FF9314037B7DEBA9303282035C0F67795417FE1;
defparam prom_inst_0.INIT_RAM_13 = 256'h93E7C8AA4C7E943D74A19B62963FF05FD33B40F809FFE6A50F33A84500CEF1E1;
defparam prom_inst_0.INIT_RAM_14 = 256'hF3A45FC1FF538383982007F9DE76DB8B71300020DB32B6C6899F14F3E1F81078;
defparam prom_inst_0.INIT_RAM_15 = 256'h1C0C0FA3F619E306818CC157BB3D886A5944763C01CBCB326DBA602FDFF20BF1;
defparam prom_inst_0.INIT_RAM_16 = 256'h8FFF5300488F936945ED426BE3783F3DBE32108665E0B81D743F37DFFF9DD96A;
defparam prom_inst_0.INIT_RAM_17 = 256'h8883822D2AC1C99140CE2FFFF8EFEA830CF000F3E2FE001842EC5EEFCB6A64EF;
defparam prom_inst_0.INIT_RAM_18 = 256'h0E4030D5379F4190F8FFC57F76E211EF97740A4FE1F4ED3327319278B2FFC06F;
defparam prom_inst_0.INIT_RAM_19 = 256'hD371A0C0FFB61099884568C7F90DFB698E364EBB574FAE5F6B77DD87FF7A03C4;
defparam prom_inst_0.INIT_RAM_1A = 256'hFDF39651B974E9B2A1877BFFC640F10820007DD5F62E643033FD8F08B9247C5D;
defparam prom_inst_0.INIT_RAM_1B = 256'h000D837FFA20BE2F827FEE3B601AD9DE399D207F6B2A3066176639FD03DEEC02;
defparam prom_inst_0.INIT_RAM_1C = 256'h38C96EE2BD004181FC00AFF813B12762E6D0337C43938D4D47F9005660030100;
defparam prom_inst_0.INIT_RAM_1D = 256'hD3F5F7386256580506497FE003008100001148368C2B0CCF8D4AF3B45FF615F4;
defparam prom_inst_0.INIT_RAM_1E = 256'hE4F217A28A43FFDFD5871F0E8A055D8EE00FB1EBE3C002FF5C33E3336B61ABB3;
defparam prom_inst_0.INIT_RAM_1F = 256'h13DF7C10F019BFBA0CB8CCCBF1F217BD0ECDF504DF85C146023FF8000010FF01;
defparam prom_inst_0.INIT_RAM_20 = 256'hE3A9DE848610A1067F761B2209F651414457466020BF02FF922673A00A370D20;
defparam prom_inst_0.INIT_RAM_21 = 256'h010E164F979EEFEFE9D2328D31F7FD20B3C552AB1A8B7203F1E125EDD26EBB01;
defparam prom_inst_0.INIT_RAM_22 = 256'h617A1E21FA5F1055DC32BED0AAA6FAF5429869CCE3DFC007E488FC0D54278202;
defparam prom_inst_0.INIT_RAM_23 = 256'h8C9A57D129E223F640BE00E6E85D036525834307DB77FB7862ABFDD07095F043;
defparam prom_inst_0.INIT_RAM_24 = 256'h400967DC5BDDC8B7813FC9A3BAF0DFCAD8B89588DFE4BD0309AAC076CCA12159;
defparam prom_inst_0.INIT_RAM_25 = 256'h4A900796828E53CC33AD3DA09B5A93A08D7D2C1D84013701F36336A3E5861F90;
defparam prom_inst_0.INIT_RAM_26 = 256'hE3CD6CFF7654485C1BFB18D56007FC100669D7D8F371DDE5A8C360DE5D3C1D3C;
defparam prom_inst_0.INIT_RAM_27 = 256'h000FFCC7E77B27A2EFA0C356590CBE4CE587F9832C18F740360F1ED119A9BF12;
defparam prom_inst_0.INIT_RAM_28 = 256'h6A1FA023314ECDE18651A201CC3BD320494047FF005387F85358D87C1DDFDC01;
defparam prom_inst_0.INIT_RAM_29 = 256'hD01741F814B06FA34160200038FFD8004EDFFFBCFCC93CFAAF9C0F7A789A0BA0;
defparam prom_inst_0.INIT_RAM_2A = 256'h87FFDF3C33875EC0F384ED94CD31D48A23F632CB633274F23C1904B080E01DA8;
defparam prom_inst_0.INIT_RAM_2B = 256'hFF953DE8C02164A8F7E829B8A72CD6D06BB17F01267BD4E57B81BE1E7FE26003;
defparam prom_inst_0.INIT_RAM_2C = 256'h7A61E7A07D65A1C8ECE09FAF9EFA101EE3083EF7F9BFE8BFC487A6F36E71C28E;
defparam prom_inst_0.INIT_RAM_2D = 256'hF3FBAB3FEEC226C220BC26448CB32DCFC8B375C904D5AAB87929CE4EA7CC4328;
defparam prom_inst_0.INIT_RAM_2E = 256'h834C7E00CCB6FC03E1DD0699C3D3AA001498D613EB1BDD58512D86094000003C;
defparam prom_inst_0.INIT_RAM_2F = 256'h26260662F03F175171381CB633300C3E7EDBF039F8FD920964FB1F100002B980;
defparam prom_inst_0.INIT_RAM_30 = 256'hA6FAFFE6EF60CC9BFCB1DD060436C24CC39FC4FDC8A816F7E4D93D2DFF98FF1E;
defparam prom_inst_0.INIT_RAM_31 = 256'h9EF2407C5467C9DB7D77F3A40E21D3FA9573283989D00905366D9CA5C200FF33;
defparam prom_inst_0.INIT_RAM_32 = 256'hDCA23E8B083C5A757B614892401FCF29E79E79DBBA23A8F42AD1576676762241;
defparam prom_inst_0.INIT_RAM_33 = 256'h96FE67D7A70C71C2CD52269C1DCDDE65BC941E53CD2D48974436234092050625;
defparam prom_inst_0.INIT_RAM_34 = 256'h0C0618625BC5ED9929D3DD3E0AE1F6F8200154172A76ABBA191DEB33804DFDFB;
defparam prom_inst_0.INIT_RAM_35 = 256'h001769A23DEFBBF040017088C3E2E587FC03845BF300BB9C2126EAD005A3E3BC;
defparam prom_inst_0.INIT_RAM_36 = 256'h61476DECC3B1A222796EEF86131FCE40F303034F3799D62D5D95CA398EE57FE6;
defparam prom_inst_0.INIT_RAM_37 = 256'hF954147ACED00ECE3C98E09BC91FF80344176B179AF0FC1580222433F8B5E3FE;
defparam prom_inst_0.INIT_RAM_38 = 256'hA8615DABF8ED9DDF6F8C26FC7DC8679CDF277B6503E500879BBAA184C9E75000;
defparam prom_inst_0.INIT_RAM_39 = 256'hAFF6F87D5AFF064B6C0038EC1F7D33F881BB0CD71C1D341FB035933E51DC2D6F;
defparam prom_inst_0.INIT_RAM_3A = 256'h6D110E0A4CCAA6798233ED1F6F5D70E4521944F6A8F9F7F86005A36F9D4F76AF;
defparam prom_inst_0.INIT_RAM_3B = 256'h2DBC25952FBFFF3A34362FEBEF7FC7E56B0F592FA44CCDBD84F89AFFFFAEEDA8;
defparam prom_inst_0.INIT_RAM_3C = 256'h69FE6D7171E66DFE280033EFEF0BE417191F3C28236D2566159B051DB7DDF76F;
defparam prom_inst_0.INIT_RAM_3D = 256'hD32B815491B9E513914C99F77FC040587E3E6C7FE843437258CCF7EE18676E0B;
defparam prom_inst_0.INIT_RAM_3E = 256'hA079046410B0ECA6133DBB8679D9A1367FE026820B92D7843804FFF7FC5898AB;
defparam prom_inst_0.INIT_RAM_3F = 256'hF8F0D320F82F601921FFFEF313F03AFDF1D35B2F6C8C1A24AABF8003FC852815;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b1;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h699065900E1B25CCC39ED3E6829971AF92EACFEF7FCF2340FEF178584621314B;
defparam prom_inst_1.INIT_RAM_01 = 256'h353245FD7DD8266E77B167A3F91116DDF4C477A44431028247F3F3A703C9D276;
defparam prom_inst_1.INIT_RAM_02 = 256'h3D062009B9FAF84EFFFF636F85DD937BBFF8F9FA630A6B1C645DCC1C6149F30A;
defparam prom_inst_1.INIT_RAM_03 = 256'hB0976EFC55F4C701816A72E82D0B921F51177F9F7504FF9DEB39F167F2BE0579;
defparam prom_inst_1.INIT_RAM_04 = 256'hA178FB4E840EBD9E7B503877C6C81B0E858DFEEE7ACD33BFFF18DAC2337A10AA;
defparam prom_inst_1.INIT_RAM_05 = 256'h5E32ADC523C58E7FFFFB1A2FD7DDC4F20CD8BB53FD40F924988799086FB7ACBE;
defparam prom_inst_1.INIT_RAM_06 = 256'h8589D23CC67F19DCB91E1F692E6A901E36F56982224F569F3B8733F11CFDD534;
defparam prom_inst_1.INIT_RAM_07 = 256'h9EF5FB0118F998F840217EA5E19300147077FDFCBC9E2CE978D9FF5DC3ACB4D4;
defparam prom_inst_1.INIT_RAM_08 = 256'h9FE4763BF70BAB487182E9B53ECC4BA3EECF9D9643B3BEED6EB259A1E2A1496B;
defparam prom_inst_1.INIT_RAM_09 = 256'hCAE0680117AB2F1D3B82846E8D1E5C0ED7FD203E3DFFFFF967FFEAF84BE408FB;
defparam prom_inst_1.INIT_RAM_0A = 256'hFF4C3F8F3FFFE61879F0423CEBCB9D91FEC9AFDE16B001A2D5FFFF836C6B6737;
defparam prom_inst_1.INIT_RAM_0B = 256'h9268F7426F008124FAA504DDA836A1CF45E0C9ADC76B90323A585C86C370857D;
defparam prom_inst_1.INIT_RAM_0C = 256'h6EB9F788F948793823BD7CDB3DB3FCFC003DE5D9F8E011F978DCAEF932430FE6;
defparam prom_inst_1.INIT_RAM_0D = 256'h13DC1F987F1AE61EFC62317CE55E7EFEA7AEA85D4F3259F4454C5A3DD4F37361;
defparam prom_inst_1.INIT_RAM_0E = 256'h2F9EBF4BA98797816821CB55D8AC307DA87A1B37B328258EB958764509483109;
defparam prom_inst_1.INIT_RAM_0F = 256'h5947C8D3E8D49602388278C0B00082809BF7E1DF8F00A76FFB63678807977361;
defparam prom_inst_1.INIT_RAM_10 = 256'hDFF67DE620E0D91CE4558049E5EC586F858F7330315FC30BC77AD0BA169AA76C;
defparam prom_inst_1.INIT_RAM_11 = 256'h75ABB68BE03DB9C4351A596AFF463E888D29A7F1E3628B1C3CFB9B08FB0543CC;
defparam prom_inst_1.INIT_RAM_12 = 256'h882FC00873A3424C3E7272464200FBF4FDFEDFF90F354BD5FE51CFE05FF5FF00;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFF58E3F548A34825DD207C63D869CA2CAB25A992C387941DB8C3A86882234;
defparam prom_inst_1.INIT_RAM_14 = 256'h0A3B92D9746DD15485AF1CC4E7B311E4782C0C5C8DCBD30441B8D2D0A3CCDEF8;
defparam prom_inst_1.INIT_RAM_15 = 256'h60086F39F5DEAC55AFABEACCB3E7FF5FDFE69138DE9F1C1336EAF221C61AC991;
defparam prom_inst_1.INIT_RAM_16 = 256'hF8324817688EC370991641F3F221E32CD658029CE5847A197DA52A597C17A20D;
defparam prom_inst_1.INIT_RAM_17 = 256'h940FDD89550B5A9AD9A4A95F06081EC72DF7C74570F3FA8F8EC5432EEAFE97F3;
defparam prom_inst_1.INIT_RAM_18 = 256'hFF4F4AFEE4EA259E55CB3FBF1429FCDBEC18EFED0032626FA5961E48B1786FF6;
defparam prom_inst_1.INIT_RAM_19 = 256'hFC737527AF0F053A884B799A87B03ECA9DFAE192B7982AC257B896E73AD2A1CC;
defparam prom_inst_1.INIT_RAM_1A = 256'h72CA59DE78D4973D921941C962AE4F0A95D78D5202FA3B146AAB7CE9BBEDF819;
defparam prom_inst_1.INIT_RAM_1B = 256'h86AC0CA16F3816069827FA73E7DE7E603FEF8A97855406362A5310E86AE982DF;
defparam prom_inst_1.INIT_RAM_1C = 256'hDBC736C10279920CDAE6DDF89B0CEBB3E51B71CA7C14B35317D1EBE6F711CA9A;
defparam prom_inst_1.INIT_RAM_1D = 256'hBA3EC5F487A1B94F36E5689A76DC3F2D3A768D7BF6AA43B5B13C54F7C1FBB8C2;
defparam prom_inst_1.INIT_RAM_1E = 256'hAB844A89CEBCF0089F927C899E9E6832B6B18FB81058049D0EAB41C24F2D2EF8;
defparam prom_inst_1.INIT_RAM_1F = 256'h36B3E47805A6220DBE87DE55E4DEC98CA45C73EBD44E21B1BD4539FD7943F9C4;
defparam prom_inst_1.INIT_RAM_20 = 256'hE9A570D31D158B6C42B88F6DE10A89AEC1CA8B50FD7C0340138FF1FF9F4F18A6;
defparam prom_inst_1.INIT_RAM_21 = 256'hD6F2361FFFD23A0B3EDFB887BD8AFF82815905EA09D230ACD28B0CD35009D980;
defparam prom_inst_1.INIT_RAM_22 = 256'h0A8438A100C736839C43C844C9A199AE0F62B9C50622BEED113F1D6C47259094;
defparam prom_inst_1.INIT_RAM_23 = 256'h71E750B740AEBABF5C035B017B891D6C496A07D3F0F082EDBFF621F600BFC079;
defparam prom_inst_1.INIT_RAM_24 = 256'h491FBE9230580466F586F5E8F02F3EC2E917284657C9761AEF16A64DE98C1299;
defparam prom_inst_1.INIT_RAM_25 = 256'h8F94447EFAEA24278D612AEDB93B06E4C4157539DC3831C6CE0FE3998C0E042D;
defparam prom_inst_1.INIT_RAM_26 = 256'h17C4EB51D9814F089BFFCF815F8E9BBCD5D0FC3254A3A6FFBF9E0E93CDA3F42F;
defparam prom_inst_1.INIT_RAM_27 = 256'hF903004F2CEDBFF79FE380ECA7711438A5F79EECA0CD9AF5209E9B8B1175E9CC;
defparam prom_inst_1.INIT_RAM_28 = 256'h3BE13B26E5C2CF616BD6A6B9F68066D6FD263F6E06405515FF3C4DEC03B049B4;
defparam prom_inst_1.INIT_RAM_29 = 256'h957CE9F0D243CA03D081B3C7FE8447BDE280BF6EDFEFF1E998A83FD4AC354F41;
defparam prom_inst_1.INIT_RAM_2A = 256'h9C0184A73DA01C66330751DEC6029D4BA69D80C0DD3449D32E014214F7A957C4;
defparam prom_inst_1.INIT_RAM_2B = 256'hFE0403FCFBD124F407D66680F1D83E26A552623449C3FC04AC96E67E30BF6EB6;
defparam prom_inst_1.INIT_RAM_2C = 256'hA69D06B0AFA73249C7BCA2BAA53F1D020EF79F89AE68FF4658D193B8222062F7;
defparam prom_inst_1.INIT_RAM_2D = 256'h9B0594EFF8F2B541E846783F9D16702144305AD3085BBA6E7BC88E6AF456BF55;
defparam prom_inst_1.INIT_RAM_2E = 256'hFB70F8EE655DBF7E16B9E504C8B97A3D9C406065410F76917DD6296CFDFD8A10;
defparam prom_inst_1.INIT_RAM_2F = 256'h09FBF8AC2D4574905B8A3CC5FF6EC42C3A647B9E39293879D56B37F9139F7983;
defparam prom_inst_1.INIT_RAM_30 = 256'h9B60BFFA778A81F44C09F604EF42457D205D232154F7D59CC82C04D0A7AD6787;
defparam prom_inst_1.INIT_RAM_31 = 256'h086871E367377FAB11952FAD4CB969DBFA164E86E2EBAEC06E48CBEF9D81B115;
defparam prom_inst_1.INIT_RAM_32 = 256'h68F0E7587620B1F5080E4AB28A52A02F017E7F7A47543537C15BCB789865FA15;
defparam prom_inst_1.INIT_RAM_33 = 256'hD9BE5F2DFEC58DEE370FEDC020586C810C443510B1F51B6D0B7F3455868063A1;
defparam prom_inst_1.INIT_RAM_34 = 256'hD2D73DCBE359C58958D19EB26060684DCD22AF10E7D09B028042C4BC448300F0;
defparam prom_inst_1.INIT_RAM_35 = 256'h1340B339C02AF5B4E357F2D17551793FF87919DC96F20709040348017394F418;
defparam prom_inst_1.INIT_RAM_36 = 256'h7EC3AFED8CC349F97799D1B8573058D2E812A03E1786B0D63384899466890729;
defparam prom_inst_1.INIT_RAM_37 = 256'h7D202987ADCE4D8A2A1DBB19A5B1A5B9468593032AD4E8876104F49208980F9E;
defparam prom_inst_1.INIT_RAM_38 = 256'hA8F47DE3890B1A98BEE16EBC77F5DF1FBD2902BA9CDB0CB6793464096E62A20B;
defparam prom_inst_1.INIT_RAM_39 = 256'h0C423B3BB8DCD10C001B1FD978B760D853293B7E045B2C3EED9DD883F6A3F561;
defparam prom_inst_1.INIT_RAM_3A = 256'hFD25D6B57CD4FE50AC9E00181A91A74F0FF5D37F006D3DBD77B795D12FFFFFE6;
defparam prom_inst_1.INIT_RAM_3B = 256'hE730BA188E9216FBE3B9F70CFFFFFB9D10CEDDDF474AFF65170DE5827608FAE1;
defparam prom_inst_1.INIT_RAM_3C = 256'h003CFED1D63F862582BF62B1390E2259AD8B122834566794118018008448F72C;
defparam prom_inst_1.INIT_RAM_3D = 256'h757FE7BDC3F85B6BC600868CDFC1F6E373FFC9C5CD61C2F55FA13E0D39E18E50;
defparam prom_inst_1.INIT_RAM_3E = 256'hFE89845387D23986C8560FB9F0FE61005ED6B1134FE059DC59B063ED7D6845B6;
defparam prom_inst_1.INIT_RAM_3F = 256'h7D86BCB60126B62FCC7EC3E5D0CEA968E061BF6FED731A2867E79241211AEE3B;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b1;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hE64F3814E33BA21859E48EC46D2E31FFBA29300FFCB2D83BD5C3EFFDBE68401F;
defparam prom_inst_2.INIT_RAM_01 = 256'hE7E7D9208BE0E9547C9FBE5E77EC4FF19DA31DD8282E29815A0DAF26F3921BC3;
defparam prom_inst_2.INIT_RAM_02 = 256'h17ECFB40EF5A37FC3ED8E30B43BEAB886351F1C0D0B82E00B9FF70017FBC3CE7;
defparam prom_inst_2.INIT_RAM_03 = 256'hECB3FFCCFA2B1F28F668C0D75C0F39F807A8177E755AF5EFB2F1F4E5C796407C;
defparam prom_inst_2.INIT_RAM_04 = 256'h324D2EEF1E5932065CF8A426D4DECB0878CEA23BB16B533365F14CD0D06B81FA;
defparam prom_inst_2.INIT_RAM_05 = 256'hD3FBC6EDA6A74FAE7F37FD55CFE7C60C03F0033C1C69EFBE8CC0780592FFCEB7;
defparam prom_inst_2.INIT_RAM_06 = 256'h23C0B11FB500FDF7EBAFFFF83FBBFCBC1F3CFD783825C1FFFFC7C66BE10768C7;
defparam prom_inst_2.INIT_RAM_07 = 256'h5A55B5121C7139FFF1F1B6FC45CF7FFBFC1A07966590946AA144B51B3373E000;
defparam prom_inst_2.INIT_RAM_08 = 256'h4481CB1B96D4CDD1EC863953F5E8C0CCF33C93EB27BF3DFAC00F3E0FFEF85220;
defparam prom_inst_2.INIT_RAM_09 = 256'hC20B986073DAF90003EDF3E7FFA2E6EEB68EDC8F9E4B9DFFCC2282E732D3E27E;
defparam prom_inst_2.INIT_RAM_0A = 256'h2C634869C8FFF61FA858F35FD463AB1D8EFAFCB4B4635E60CE1305F3EF3CC00B;
defparam prom_inst_2.INIT_RAM_0B = 256'h819A58E9FEDFA8AAA934D37A1F3BF360C96EA603977D10C0059EF7B9E123AC58;
defparam prom_inst_2.INIT_RAM_0C = 256'h1BC980FDDF8400018C9E6FF85656C49BC8AE3073FFFD9FF2160CEC0722E586AA;
defparam prom_inst_2.INIT_RAM_0D = 256'h4A0AA2F927FBEFE8655321F3FE764BBF9B1CCABC0D8AF3C3AAD3610FDDFFD80F;
defparam prom_inst_2.INIT_RAM_0E = 256'h8DC523E490A2A89A4D607C0CFC6006B2E4008DF1C07CE6AD966BFF1E74AF01A7;
defparam prom_inst_2.INIT_RAM_0F = 256'h80237C780F789FD11F79C062AAC70CE902EBA84D9F7C583458572ECF5B0499E0;
defparam prom_inst_2.INIT_RAM_10 = 256'h1363FEE07FDF28DFDB0BC7444040980B70B05AD0BCD47A5520C203302C0DAEBA;
defparam prom_inst_2.INIT_RAM_11 = 256'h8FFBC4A523FB7B581008070043FE838063F7FFFFF181FE04F9F9806ECDFE7F36;
defparam prom_inst_2.INIT_RAM_12 = 256'h85B55AE6A01BA94EFD80EFB965BD9222707BBEF7A72BECD79C2CD890177E688F;
defparam prom_inst_2.INIT_RAM_13 = 256'h7EFFBBE9CA07F9C4CD856CA9C780637CEFA6C74CD382DD1A00FC9000F2E0E001;
defparam prom_inst_2.INIT_RAM_14 = 256'h2975F32988F742983F2B003FB84180016CF56B6F263553BF6223F1DF00B452EE;
defparam prom_inst_2.INIT_RAM_15 = 256'h7F17BAF4C2E3FB86017FCE42B71AC27396FF6696E1AB016030334A71E40020C7;
defparam prom_inst_2.INIT_RAM_16 = 256'hFFE7663C1355C8B0007EF9DA5F023C475D62F005ED1880D1B0A30FDF2E021800;
defparam prom_inst_2.INIT_RAM_17 = 256'h7110D92F5820072235B33BB9F0070C58DC935085FAC04021C065790F58180CF1;
defparam prom_inst_2.INIT_RAM_18 = 256'h05D8C17FD0100802028EEFDD6E8438FFE7DB2F11D553B4817D99A1281044DF90;
defparam prom_inst_2.INIT_RAM_19 = 256'hFEF6D7B12BDC103219F1D784A03699F928700A10098EBD7390CEBBE3843C9D25;
defparam prom_inst_2.INIT_RAM_1A = 256'h3EAFC36112C00B4E0E4156B2FB5BE13E3C0003E65B001BB4347E7760E1A5AF1B;
defparam prom_inst_2.INIT_RAM_1B = 256'h8000F9F7B806ED01DE21A3CFA4EBC7693BB7EC2317511F2CFF77E39B5320FF91;
defparam prom_inst_2.INIT_RAM_1C = 256'hFECE6C2A5441D371D438DD0C8F3FEC833B10B8A05601CB839C50306EB6FEDB37;
defparam prom_inst_2.INIT_RAM_1D = 256'h7B6E0E2C00C469D0011CB8A3800C0AFC03EE96107137A1FF7CE6BFFAB6CB9BFD;
defparam prom_inst_2.INIT_RAM_1E = 256'h0667C5183CFF00C2B1051D84DA7EFCD97DC252F11C864FE880FC9D1F264C0E0C;
defparam prom_inst_2.INIT_RAM_1F = 256'h71A1F4C081037F4028F8741C3448B12E11200364F18C000019B1860012804F80;
defparam prom_inst_2.INIT_RAM_20 = 256'h480219FFE303D78A9E518007A0D2E80D4192248EDF001C1F2AAEF736DE5EB64B;
defparam prom_inst_2.INIT_RAM_21 = 256'hCF85DDAFFC21CB4CFF7C68FF9FD7FFF85C7630A6016F980E2CFD331C53B31464;
defparam prom_inst_2.INIT_RAM_22 = 256'h94BD1307D0757E126783EA0EDEB3D98A04AA4FAD7C07AF4FC07FFEE2193BA17D;
defparam prom_inst_2.INIT_RAM_23 = 256'hCE077F13FFE4439787E962871ED957D9E055EBFFF92272F3110047B1C8FBCA3F;
defparam prom_inst_2.INIT_RAM_24 = 256'h577AE67C075D6FB6080185F99ECE8E539F631E0300E083E134725A9DFAC38E03;
defparam prom_inst_2.INIT_RAM_25 = 256'h58DC05C05E23B0FF0059A154ED33E0D581DFE7FEDE03C5F80D5745047F41EFF0;
defparam prom_inst_2.INIT_RAM_26 = 256'hEDD1AFF1A797A02000CFDDB6940B94143DFFD7F03C940257884D07733FFF2CDF;
defparam prom_inst_2.INIT_RAM_27 = 256'h78FACD00E61142B210BB73903CCAAF064DCBCCF31883EC234248E78D5DCB6D68;
defparam prom_inst_2.INIT_RAM_28 = 256'hF092C3C8F30708604AF56AB173350A37756995B903F850BAFBC05D924E91F249;
defparam prom_inst_2.INIT_RAM_29 = 256'h2E052464A40E2C854FC83F2520AD126F6F9E43434160F170299B379F770BC051;
defparam prom_inst_2.INIT_RAM_2A = 256'hADCCB0B27B0AF4E1B4CE7F36120AC60A81DA324A933864784261611FE88687F9;
defparam prom_inst_2.INIT_RAM_2B = 256'hCBE5F024D8537BE3EB954EE00A12FFD5AB61E06EB670787EC815D8A881231737;
defparam prom_inst_2.INIT_RAM_2C = 256'hC8F81C22B534DF820E2DD61228BE9DCBB30743A6450AD9F553D0FCBC14114948;
defparam prom_inst_2.INIT_RAM_2D = 256'h80DEB41ECBC9CC7EE7F080388035FBBEA01C8B329B3C1174DCD3F85AA87FCF0B;
defparam prom_inst_2.INIT_RAM_2E = 256'h29E0439603E57EFB706EB979CF071FE0FBF9D9877108803098DC758B26236D1F;
defparam prom_inst_2.INIT_RAM_2F = 256'hFCE0EB6802E00015D67640DD7925F3E0F30DE506BF89AE6F842A1D4E97E2A790;
defparam prom_inst_2.INIT_RAM_30 = 256'h468EEDE3204F5DF6D4F8CC45EABC9E300011221F770E49C43749B51702C362FF;
defparam prom_inst_2.INIT_RAM_31 = 256'h3780CA9F944F8F1F199AD3C1FB7E6BD8EA53981F42027B9540C01E0062FEFB0F;
defparam prom_inst_2.INIT_RAM_32 = 256'hE68007C8410DB83FEF9E003DB334277EE29D4E8F6EF60A123CE4522E2E841514;
defparam prom_inst_2.INIT_RAM_33 = 256'h8CCDC3DBBF92C4B771104BAF00E1A01CA5EAA13DAECF47F00FDADE5A2ADFFCBD;
defparam prom_inst_2.INIT_RAM_34 = 256'hB92C96161271FE25F86EAB10FB98D49B2639F220B01ACFDBE643B361CE041069;
defparam prom_inst_2.INIT_RAM_35 = 256'h88EFF366A3B79FFF9E85BEB7BC1347F6A906D8987C60515FD452E0904718CB5D;
defparam prom_inst_2.INIT_RAM_36 = 256'h75B90739C11AEDD2B070600288003C21312D7E2CC61D713F0FDF5BB778FC08F9;
defparam prom_inst_2.INIT_RAM_37 = 256'h14F1D791A5FBEE00713E93D0D17E0643057C6340397FDFF870A2CFFD32E4CFE5;
defparam prom_inst_2.INIT_RAM_38 = 256'h6F9A57CE9FF7F81E1094FE4CB60D6010D3464EB38EBF4C959B90566218D4178D;
defparam prom_inst_2.INIT_RAM_39 = 256'h09804FE3AE99E458C19D1886270AEB9459F38C087E7B0C12EA58F17FD67F8841;
defparam prom_inst_2.INIT_RAM_3A = 256'hBB8EE0047648384AA8F8B64BBBC042FFFE7AA60DAFFF07F1EA4E0D7DCB43A65A;
defparam prom_inst_2.INIT_RAM_3B = 256'h03DF816DEDDDD91FD000F754D7C9A59E879979CF3F22C00122F7E7FF61673E01;
defparam prom_inst_2.INIT_RAM_3C = 256'hFE5733EF05B5A39D91FA1FC5D67A67ACB3C809B6BA60F58609DC3E8FF60025FC;
defparam prom_inst_2.INIT_RAM_3D = 256'hFC0001009DBCA880C74E089FA18FF3BD4F1D3EFCDFFF2DC6433FD8564EEA09A1;
defparam prom_inst_2.INIT_RAM_3E = 256'h2DE1A17F7FDBBAFB3FF432DBE7DF1485F60F18C2008666ED6A03BD6335337B71;
defparam prom_inst_2.INIT_RAM_3F = 256'h4B2F1F963DF833B7BFCD1162749DA67810C3900CF121A3763F001BE01BEF3504;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b1;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h528403D95368F72840017844FBD1A6F478713FD7F6B20EFFFC0E6679D5728183;
defparam prom_inst_3.INIT_RAM_01 = 256'h00806A9EF1766C7DB3F7A089BBDECA70640312A6EE2973F3F0B259DA8A6B9802;
defparam prom_inst_3.INIT_RAM_02 = 256'h7D9DA9B687FFFFFFF96FE05847CF8D00260FDC67EFC71E40007F810071B699FE;
defparam prom_inst_3.INIT_RAM_03 = 256'h2FA724FEFE3F861857FA1000241FFB7997667C122D1ECFB7CEA94B386CD95730;
defparam prom_inst_3.INIT_RAM_04 = 256'h41A706A093702DFB1B8B132B3E90DCC82E13EEE8FFEFC2877BA50D74DF8E18CA;
defparam prom_inst_3.INIT_RAM_05 = 256'h40FE9C39BD98902EA9E369A3E206520BE79F238E2D600011FFE40819D28FB684;
defparam prom_inst_3.INIT_RAM_06 = 256'h94F1EE10BFBC005F5B2028CCFEEA7FB006010586EBFC2FE99105AD0BBDC64D08;
defparam prom_inst_3.INIT_RAM_07 = 256'h027F73A8FE77F836B4859C975D8F07FFAAA0A17C6C11B06616DAE9E73F278385;
defparam prom_inst_3.INIT_RAM_08 = 256'hC928373B473F93A1139A7E562C70C352D02223EB0B7E1FFF7A7BC5C46BFFFC47;
defparam prom_inst_3.INIT_RAM_09 = 256'h075262FEA0165FF432D7C8637FB691829C72E1780FEE1442C44A67E27332CE4C;
defparam prom_inst_3.INIT_RAM_0A = 256'hA9B8210CFE1F1E3CA7055F103EBB4FDDE206021BEABD9EF2D5E6E7FDE6F46FCA;
defparam prom_inst_3.INIT_RAM_0B = 256'h438C47CBB5A56CA21E7FF9FFFBA582A09877FBFE0D231C04354850637FEF9C7F;
defparam prom_inst_3.INIT_RAM_0C = 256'h63FEFFE4CAC7010C47580ED8637F19EDD574C37F81CE0F05A682D73499EE561F;
defparam prom_inst_3.INIT_RAM_0D = 256'h0828F0AE3227BA583BEF9EC278CD87C8E493C2E14A602FC63FFC5FBE253947DA;
defparam prom_inst_3.INIT_RAM_0E = 256'h6049F80E37D7A1EE47FE3B3E4C91477C1DF7FF80483A26D92BCFF7F7FFE9FA1F;
defparam prom_inst_3.INIT_RAM_0F = 256'h6FA7E000D7832C8AC8FF839D2D188E5F2D47CBF1FD6865D0EDE1130F7FE18596;
defparam prom_inst_3.INIT_RAM_10 = 256'h5EF224C8129177DB4153C8639646E41565BD5C9E9DD92FE9BFB18A3CEED35233;
defparam prom_inst_3.INIT_RAM_11 = 256'h22B27700D6CBFDEFEB6201C7B9DAFDBB9FF801CBE3F8FF9F7F8E9F337EA609C8;
defparam prom_inst_3.INIT_RAM_12 = 256'h65828C3439D6DBA6AFFAFDFE8E6D3C1EDC80F3CB6F15F208F49E766689A10529;
defparam prom_inst_3.INIT_RAM_13 = 256'h38400D829613FECEDF267EBCD80FC30AEE211C09F1FBF7FE6637FF4DDE1A65DF;
defparam prom_inst_3.INIT_RAM_14 = 256'h2404AF447F67FFB6DF28CBE20EE967DAD8C00E0EBA577A9DF8FF7FED641FFBFE;
defparam prom_inst_3.INIT_RAM_15 = 256'h7E01EB0FA3D8A3FF8AFFF96E5BFE288104CEBAF0132EBF85E4DC2F093A7B1093;
defparam prom_inst_3.INIT_RAM_16 = 256'h2979E1B231FB6FCB369501EC4C5EF42ADB3C3291FFBFDC52713E11CFB8F41EBF;
defparam prom_inst_3.INIT_RAM_17 = 256'h7B0CE38E6E681DBEF72BA84FB1F413F7E83EF72F649E6CBFBF7FE9083DE28274;
defparam prom_inst_3.INIT_RAM_18 = 256'h037C8B0ADDFD2BEFC7C46F3F76A0151C936524F6BED568EBDE307810BF31A0D2;
defparam prom_inst_3.INIT_RAM_19 = 256'h16A641E1956A2877E41FEB0E932AD5A3333F7A1BF60422FDC689D3ED7C1CFDFE;
defparam prom_inst_3.INIT_RAM_1A = 256'h940AC56212ED4EC109A88618417E5F41DB0B3FF51C0A7E7B88CC87FB460BC628;
defparam prom_inst_3.INIT_RAM_1B = 256'h3492376501F9CD472980CB33010360919CE3B624CE22E8E824647903CC67A241;
defparam prom_inst_3.INIT_RAM_1C = 256'hC5F3F920F32803ABAA485207F022E4695181A61FFC3D23C7991F91A027F4FF30;
defparam prom_inst_3.INIT_RAM_1D = 256'h611701A4FC4887AE47986110797FF4023B63CA187F7736ECB404C8000158D772;
defparam prom_inst_3.INIT_RAM_1E = 256'hE7737BC0FECD57960019868F805EA5B83E53A8D4FB18E0901ABB1FBA19A96854;
defparam prom_inst_3.INIT_RAM_1F = 256'h55F9F1F77844EAC285C62EAF781339F96070099A81F468E186016001D6CFD47F;
defparam prom_inst_3.INIT_RAM_20 = 256'h9BA35D43B120397FE6164670BDFD0B3A2E19BA6742B2FA030D66B3800E7F2DC9;
defparam prom_inst_3.INIT_RAM_21 = 256'hD748AFDD6EDB8FCD012FAE02C275F2E3357E817E106DD5F844FFE8557BE96639;
defparam prom_inst_3.INIT_RAM_22 = 256'h89C4378A2238A05B9CF0902BFE2FF19DE3A260DB15579FD8595F6C0E943800B9;
defparam prom_inst_3.INIT_RAM_23 = 256'h8A0CFDDD0D4BE68FFFFFFCF0088261F5CB274D6B67857CDABC96B8724368B78B;
defparam prom_inst_3.INIT_RAM_24 = 256'h96F5EDBA1D6CF74F7FCE1A10B0DBF00FF082022C06070722AC7318299BBBF7FA;
defparam prom_inst_3.INIT_RAM_25 = 256'h28808A8F6A2A8E9C93A697A7779DFABDDF30C57D737DFB9FEFC7C3EBDF175827;
defparam prom_inst_3.INIT_RAM_26 = 256'hF87E0FD49DA1523F8A23450B9979847F84FFCB65302610C14987C2568A67C3CC;
defparam prom_inst_3.INIT_RAM_27 = 256'hD506063C2DF501A453C6FC98665F00DE34E1970BF6A0E25B17786DF3D97D2E59;
defparam prom_inst_3.INIT_RAM_28 = 256'h10FB72BFB9C30A5A7FAFF3CB4818E3C1464421567FFF138A0A3B09864271DDC3;
defparam prom_inst_3.INIT_RAM_29 = 256'hDB08459EE1C49B722D0021EED179005F01208F0BF280110B08E13991A5E7C1A8;
defparam prom_inst_3.INIT_RAM_2A = 256'hEC22E620115823FFABF11A4FFE3C6E1A60C3EAADE53D124CD8FEF6CD87BD30EE;
defparam prom_inst_3.INIT_RAM_2B = 256'h72A149B2E12CBD2AB97FEFE7973FCEB83479E0018AF9509E404A40A7BE107173;
defparam prom_inst_3.INIT_RAM_2C = 256'h4D11078CDFB9EBBD84B40F2F9E9CD20347B4612C468E9FE70BE7C0C817E62E8B;
defparam prom_inst_3.INIT_RAM_2D = 256'h828F013C4BF983DA308337C5FE23A22B0678D4244B8D05869FDDE1E987CC16DD;
defparam prom_inst_3.INIT_RAM_2E = 256'h13993434695E5468318878E40B9DCB8B5F0601F900B19531A7E1DECD290CFE0B;
defparam prom_inst_3.INIT_RAM_2F = 256'h87C7BE25088B9A8C1DA9131B3EDADF84C1CBFA5A5275881F4E3218F04B9AA4EE;
defparam prom_inst_3.INIT_RAM_30 = 256'h32FEC695057230EC7046895E77181F57CFC61D695CA6357820D0F51B680BDEEF;
defparam prom_inst_3.INIT_RAM_31 = 256'hAB7C53A4F22B3E0830C50B192BF78DE9F1EF89423AF4C16A0B5DA517D6FC29F0;
defparam prom_inst_3.INIT_RAM_32 = 256'hB77C66CB9D9BD64E08C50E58EDA6CC1F4C981007AA8918482D669CDC3C557A35;
defparam prom_inst_3.INIT_RAM_33 = 256'h566700440B78D08987313CB47A83B40E4CEECF7E777C219D01029531E4EB7CD3;
defparam prom_inst_3.INIT_RAM_34 = 256'h357ED1AA7E7B77B52B225B450C6FFFC6816193E1C7078F6409F9A5E586E9C297;
defparam prom_inst_3.INIT_RAM_35 = 256'hD9377EA4B618443E6DF17965259F9535104429634A7FE8BEAA7E5FB5A844953F;
defparam prom_inst_3.INIT_RAM_36 = 256'h8E19C79005D57B94B39DA8B2E8D9137FDAE0DF19DEDB6B67CB9A5C431A63EFB9;
defparam prom_inst_3.INIT_RAM_37 = 256'h18009FA867E35C68A101B97873185866AA149A12A80BDABB97FD9060C736352C;
defparam prom_inst_3.INIT_RAM_38 = 256'h5CFBAA59D097F01BE81B1830FE014F6D818D8662E9B802E2F647E7548AB3758E;
defparam prom_inst_3.INIT_RAM_39 = 256'hD02A64675D024636D5AE79962236EB40A896EA3C71481E2607DE561D58F7E123;
defparam prom_inst_3.INIT_RAM_3A = 256'hC84F7EF8226F614941042729982864D7617F9B2FA089BE7DF87D743942111841;
defparam prom_inst_3.INIT_RAM_3B = 256'h9D6DA9F59AB77B0E12583F53568119D90948710322B04DFA9F88E7A4B2758581;
defparam prom_inst_3.INIT_RAM_3C = 256'h13AE9368C29B6EFD7D603FE85BB3DF024EF74DFF11847D8309C7401045DDD69E;
defparam prom_inst_3.INIT_RAM_3D = 256'hBDCA59446EDD7FCE71480450ECA82A14DD1D6AA5CBC4C3E4A60C20C74B8C77C2;
defparam prom_inst_3.INIT_RAM_3E = 256'h1AB9DD32B60FE6C4F3E01814350918B1EBBAD3322621FA00E18B1B86C37720C3;
defparam prom_inst_3.INIT_RAM_3F = 256'h74E42DC1865F3CBA3661D22EE300FE1B8060D04485BC9715D0727F07646EE2C7;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b1;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h0005007931E9FEBF9FFDFFDFEFFFBFFFFFFF679FFFAE00004004DEEFFF7C0BC0;
defparam prom_inst_4.INIT_RAM_01 = 256'hBFFFFFEFEC0000105EAFD8295CC4E86B7A54404000C9425FFC801397FB800000;
defparam prom_inst_4.INIT_RAM_02 = 256'h97CCC8832FF2F73D2014FFF620000810C4B330403E7EFBDF766FFDFF87DBEFFF;
defparam prom_inst_4.INIT_RAM_03 = 256'hBFF821597FFFFFFF7FDFFCFFBA7FE7FFDC6D9FF73C70000006AFFF9BFC3FA1E5;
defparam prom_inst_4.INIT_RAM_04 = 256'hE7DDD7FF542101800BA69FFE616876E4C0EF0204434EFB8804BFFE100000E07F;
defparam prom_inst_4.INIT_RAM_05 = 256'h8011302B5D73C082EFFAC0000058A3FB3F8001397DFFF9FFF7FFC819F61D8007;
defparam prom_inst_4.INIT_RAM_06 = 256'hE000184EF7FE79FFFF300210006001999A76FFF90850200171D9FFE077FFBA01;
defparam prom_inst_4.INIT_RAM_07 = 256'hE0FCFF4C8E04412005E7BC03BFFC8078004C3CDFFC0000BFFED11E000228FEFF;
defparam prom_inst_4.INIT_RAM_08 = 256'h0009FFDD20005FBE400000196E3F7F9F01021B79DFFFFF4C0209101108032B43;
defparam prom_inst_4.INIT_RAM_09 = 256'hC900637FB41E8600000040400B664A2D02CFFB3C000800007967EC6FDB0A0092;
defparam prom_inst_4.INIT_RAM_0A = 256'hBFFFFF00000000066DE01FF712003D0043DFCF0C202FB20880004BB7F7CFDFB0;
defparam prom_inst_4.INIT_RAM_0B = 256'hDFF1C3042FEF42400017CAE20FF7EC005818FFE807A0800008205402C86A8860;
defparam prom_inst_4.INIT_RAM_0C = 256'h01FF8696003008200445001049C0027FFFD7EF682008855EFB8BD8C320801869;
defparam prom_inst_4.INIT_RAM_0D = 256'hCB3DDB580026532BD8DFC51800020DAFE74C348EEF74000008F8D4EBBFF30000;
defparam prom_inst_4.INIT_RAM_0E = 256'hD80623FBFB000006F42FDC2FCD0108007FE020800C0180100880001A800037FD;
defparam prom_inst_4.INIT_RAM_0F = 256'hFE068000000200000000184E081FFFBF5BFF1001001C0BCA87515C624C622FEF;
defparam prom_inst_4.INIT_RAM_10 = 256'hFFDD20000A6C3797C03014E179FFB6E2108FF6F340000A98F5CBFBD3C000241F;
defparam prom_inst_4.INIT_RAM_11 = 256'h007EFD008006102EA4BFE001100539F786441C000000003000038AFF0DFCF7FE;
defparam prom_inst_4.INIT_RAM_12 = 256'h910300000000080000E22DC1FFFFFEBFE84820028303D460002A080A697D7FC0;
defparam prom_inst_4.INIT_RAM_13 = 256'h640000080475F0000100240FFEFFC0202FBB40400FFA4DB1DEC2A04100CFFBE1;
defparam prom_inst_4.INIT_RAM_14 = 256'hFFA4000BBDEA27FCDCE007F9FE7FDB837040000000151090009D1C73FFFFEF9B;
defparam prom_inst_4.INIT_RAM_15 = 256'h10000C50004C000001844F59FFEFFED787B3847805FBC10812001FFF5FF0040E;
defparam prom_inst_4.INIT_RAM_16 = 256'h540001003E04809032029DEBE000C0DFFE000DFBAD55371F973FF7DFFFF9F962;
defparam prom_inst_4.INIT_RAM_17 = 256'h800076CD0D93CD997BFFFFFFFEEFF88800F000000000008042EC5FEEFFEFCF20;
defparam prom_inst_4.INIT_RAM_18 = 256'h0240018100000000F0FFFDDDFBEFFE184880000E800042C898C7727880003FEF;
defparam prom_inst_4.INIT_RAM_19 = 256'h200C00C100019627FFBD788406F3FB6804FFFE07BEFD8CABBFFFFFEFFF7A0000;
defparam prom_inst_4.INIT_RAM_1A = 256'h09FFBB1621E74947FFEF87FFE6C00000800068400100602233FFF9BF7EBF8322;
defparam prom_inst_4.INIT_RAM_1B = 256'h0000800001803D3FDAEFFFFDFFE72221888030804045DF9DFF0F11027FAEC400;
defparam prom_inst_4.INIT_RAM_1C = 256'h0048101402BFBF7FDE000007FBF127897ABC6FBD4923F13DBF87FFBE60200800;
defparam prom_inst_4.INIT_RAM_1D = 256'h45F0677CD27B9BFAFFB7FFE00000000101010000000B0EFFCEFFAE5F7D8DEA03;
defparam prom_inst_4.INIT_RAM_1E = 256'hC0A0000002C3FFDFDFEFCBD7FFFAA240116242059C3FFFFF580014DFEB628CC1;
defparam prom_inst_4.INIT_RAM_1F = 256'h00D1821F0FFFFFBA000537FBF03FE150B5242380DBFF3FBFFDFFF8000000FF01;
defparam prom_inst_4.INIT_RAM_20 = 256'h869E008026EF1EFFFF7618000BCCE5400055002020FFAFFFF7FBFFFFFD98F10C;
defparam prom_inst_4.INIT_RAM_21 = 256'h0100004F97DFFFFDFFBF7DF8CF0012265C22AD44F7FF7220000FCFFCAFE8799A;
defparam prom_inst_4.INIT_RAM_22 = 256'h048461DCE7FF100023EFBF87FF73686A9D5AF2098421BFFFF48100059A2D8600;
defparam prom_inst_4.INIT_RAM_23 = 256'hFB6434A5061BDDF640000129222C000025010307EBFFFBFFFFFFBE2FC7608234;
defparam prom_inst_4.INIT_RAM_24 = 256'h40016FDFDBEFFFFE7BFEFFDE01088090275F6A7FDFE09070F6FBF7EFF56C9EB7;
defparam prom_inst_4.INIT_RAM_25 = 256'h95FFFF9702860833F3E7DDA54665EEE7C76090001BFEFF400C829BC42D804040;
defparam prom_inst_4.INIT_RAM_26 = 256'h28F13C9889AE4803E304102F601000100269F7F9FBFDFFEFFF77FFA0220002CB;
defparam prom_inst_4.INIT_RAM_27 = 256'h000FFDFFD37B3FE7D5DF7C89A20A31B73AFDFBA0000208BCC9B77D66569E4090;
defparam prom_inst_4.INIT_RAM_28 = 256'hBEFF80030091F3EADFD1D89872084FAB5C0000009FF0002015F4C63A00200400;
defparam prom_inst_4.INIT_RAM_29 = 256'h74B74007FC819024A16D8F60060000000EDFFBBCF8D97FFFFCFFD081A20175C7;
defparam prom_inst_4.INIT_RAM_2A = 256'h87FFFF3F32DFFFFDCF79124B224E7BF3FFFE200010CDBF22DDF41E5595FF2AF3;
defparam prom_inst_4.INIT_RAM_2B = 256'hFF9404073FDF4678BD81D7D1D00BB9B91FE1007D20041E2EBBE4C60180000003;
defparam prom_inst_4.INIT_RAM_2C = 256'hFE201FA002070E0C2CCB90506100001EEFFE7FF7B9FFD3FF5F78110C819BFFFE;
defparam prom_inst_4.INIT_RAM_2D = 256'hF3FFFFBFEEDFFFFFDB43DFB3735FFDCE90800017FBE72451B67ABDE9082A5FA7;
defparam prom_inst_4.INIT_RAM_2E = 256'h004000FF31589C000DF7EB40328FADFFD487D60043B2E8B9C89C19F40000003C;
defparam prom_inst_4.INIT_RAM_2F = 256'h01E60204E2B0CE770B06E34000000C3E3FDBDDFBF1FDFFF6930000EFFFFFF988;
defparam prom_inst_4.INIT_RAM_30 = 256'hB7FEFFEEFFFDF3E4030E22F9FFF6E80000003BCE00A6C109BBD3F41F86B980FE;
defparam prom_inst_4.INIT_RAM_31 = 256'h800DBF95E924A68B3CA80942BFA02FFA7D40003DDF6FE1A2709362000000BF3F;
defparam prom_inst_4.INIT_RAM_32 = 256'hD0203F3027F4EDAD04BC5880001FCFFFE6BEFBDFFFFE770A3426AD96F2742000;
defparam prom_inst_4.INIT_RAM_33 = 256'h9EFE7FFFF3FB8E0D32AFD9BC19488400436BE85DFE90B1CA338E6ABE8E02FE1F;
defparam prom_inst_4.INIT_RAM_34 = 256'hF7F91AE22018CE74D42C33EDFA1FCBF800016261FAA63985E61DEA01004DFFFB;
defparam prom_inst_4.INIT_RAM_35 = 256'h00114787044CF81788001080C3EEF597FCFFFEFFBBF744037FFBFBD001A00002;
defparam prom_inst_4.INIT_RAM_36 = 256'h6167FDDFFC8654DD9EEFE984000051BF4C9328EC0867337E48B51F0781E2FFC0;
defparam prom_inst_4.INIT_RAM_37 = 256'h0DD6296F316E39E72702607838FFF00047BF4F9F5BAE03E580062433F8BFE3FE;
defparam prom_inst_4.INIT_RAM_38 = 256'hCA1B5C5E77226026020026DCFDFBF7FCDF7FBBFE9498FF7E7BFAA1000000AFFF;
defparam prom_inst_4.INIT_RAM_39 = 256'hFBFEFFC2A401C7BFEC00009000808C030C75032EFCFADB02186F8F0E2DDC284F;
defparam prom_inst_4.INIT_RAM_3A = 256'h9A6C75D7DEE0214685F1E302FF5D73F93FDFC15FD80000002001A37FFF4FFFAF;
defparam prom_inst_4.INIT_RAM_3B = 256'h4B007C93004000002037FFEFE77FA7E7693FF0C04BBFBF7F84589800005101FA;
defparam prom_inst_4.INIT_RAM_3C = 256'hFDEDD0DA9FFEEDFE2000041010F0314A156FD3BBBFC0C4AB8F78C2FFFFDDF84D;
defparam prom_inst_4.INIT_RAM_3D = 256'hE78C3ED4C02C780B4F3C67FFFFFF84684504FC30071C800058CCFFFE19E76E1B;
defparam prom_inst_4.INIT_RAM_3E = 256'hAC864C0BA7000026333FFF9E79D9E3FF7787D97DFFFAD784300000080059670D;
defparam prom_inst_4.INIT_RAM_3F = 256'hE38D2CDDFB2DE0912000010C12DBA9628F28B0745E8D391387807FFC03591E0C;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b1;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h3C6A18003E075343C04116BC4010B7226CEFC01080B08B40FE75F87E4423310F;
defparam prom_inst_5.INIT_RAM_01 = 256'h3510BA02000037FEFFBFE7E3F93D77F49B3F29EFC531028000800427E1EF3FDA;
defparam prom_inst_5.INIT_RAM_02 = 256'h8FF9B6E9B9C8F84000000370A3B34292426C35E52D46D8FC0017D703C043441A;
defparam prom_inst_5.INIT_RAM_03 = 256'h617E4CF70DAC3F01F24A4BCC288B82CDD70080400004FF9FEB79F167BEFD6F00;
defparam prom_inst_5.INIT_RAM_04 = 256'hE0870400848EBDFFFFF03877DFD7C6617FFFFEEE784D30000000D8082CE9F1BB;
defparam prom_inst_5.INIT_RAM_05 = 256'hBFF6FDC523C78E0001FC0704457AD00162AD39D92B6FF1C9E14D79FE3954BD08;
defparam prom_inst_5.INIT_RAM_06 = 256'hA0B81149C9FFE9BF159149E692637C6601021202236F779F7B873FF9FFB26BDF;
defparam prom_inst_5.INIT_RAM_07 = 256'h610A00015FFFDEFE40807EFFFC6CFFFFFCFFFDFEFC9E00017F13EE56DBF55C26;
defparam prom_inst_5.INIT_RAM_08 = 256'h9FE4767BD7000B4B807F10C2B2C026329FAECD71BEC66026D324C2CB1AFFCBE0;
defparam prom_inst_5.INIT_RAM_09 = 256'hD924D87EC37CE1025066EE5312C7BC112800003FFDFFFFF967FFDFFF041F777B;
defparam prom_inst_5.INIT_RAM_0A = 256'h000C3FFFFFFFE6187FFFFFC3167F6FDBFEFFFFFE1E8001433E1EC284F8992077;
defparam prom_inst_5.INIT_RAM_0B = 256'h97FFFF4BE100F9DB01ADCD2D74DB03FA29BF864E7C7CD9D1C984079B57B78002;
defparam prom_inst_5.INIT_RAM_0C = 256'h19A006A18343B0405A2A479C1D702102002CFFFEF8E011F978DED806EDBDFFE6;
defparam prom_inst_5.INIT_RAM_0D = 256'h13BFDF9E7F1AED1FFF76018B7FFF7EFEFE7EE3654F7C6E65B86BEC864EB2B66B;
defparam prom_inst_5.INIT_RAM_0E = 256'hF61C544FB21B8D161A5E14BF8890BE0C6801782EA3EB262FB4734BB34F400D00;
defparam prom_inst_5.INIT_RAM_0F = 256'h21B4E420053940A7BD157EF6700000009FF7FFDF9F78A7EFFCAC1F7FFFFFFBFF;
defparam prom_inst_5.INIT_RAM_10 = 256'hDFFFFDE7A0F8DDFF03286FEFFFFFDFC225D0E27DC62BB8F4A6A430021CDD671C;
defparam prom_inst_5.INIT_RAM_11 = 256'h56E311F1ABB9C785F13721419A378680CB8379811E6147BABED8DB47FB0003DF;
defparam prom_inst_5.INIT_RAM_12 = 256'h90F5BFE52CCE3E80B1762E3E4200FFF4FFFEFFF90F375F3000AFF7FFFFBB6376;
defparam prom_inst_5.INIT_RAM_13 = 256'hFFFFF3847F7DFC032FFFE5EFBC5BC21BE0EB8C68982BCD414A68A8179BC1A021;
defparam prom_inst_5.INIT_RAM_14 = 256'h086C1D015DFDC9C54D6103C7B4701B1A219C0F7E7BB7F1D8A86D49D023CFDEFE;
defparam prom_inst_5.INIT_RAM_15 = 256'hDC007462F0A75FFD6023D4CCF3F7FFFFFFE69118FEF202CCFDFF7FFE4731C8A7;
defparam prom_inst_5.INIT_RAM_16 = 256'hF932481FDFC81C9FFEFFFE35ABC3F42FCA1E78F6353FAA5BEB7DBB930C050E65;
defparam prom_inst_5.INIT_RAM_17 = 256'h450903851B034E8E7F6AED43073976CF12067D7C38395D1F2B92933EFFFCDFF3;
defparam prom_inst_5.INIT_RAM_18 = 256'h006FF8F7CA0AC8F1BF61FFFF35F9FCFEEFBCEFFFF0443FDFDFFFD5159FFC7FFA;
defparam prom_inst_5.INIT_RAM_19 = 256'h707BFFC991F9FBDDF7B37E57086580731E2D8793D89BF315D7895DE7CB37F783;
defparam prom_inst_5.INIT_RAM_1A = 256'h3C9AF232A73D889A397E3BF70DC7C8F427E07562E01869CFEE1FFCFBFBFFF859;
defparam prom_inst_5.INIT_RAM_1B = 256'hB331C4310C45D3FD80FFFEF7FEDE7E603FEFF0B47AF9BF8DDC4CCEC9F8E10198;
defparam prom_inst_5.INIT_RAM_1C = 256'hF9DFF02EFF17FDF752FDF9BEBCB0CDC9C0C89E233ED6046E5E8FF25D41703D60;
defparam prom_inst_5.INIT_RAM_1D = 256'hA9820127A792E7D571FE1F7BCE0BC03DDCC08B638D1D3034AFBEDBF7E1FBBA82;
defparam prom_inst_5.INIT_RAM_1E = 256'h9E353E30B4C00D0BFFBBFC99DE975030F700001FFFA7FD7267B79A6B8C36429C;
defparam prom_inst_5.INIT_RAM_1F = 256'hCAE01B8BF7F9DE0D4BE46628396B58C255A5FFECE2336A087B89779302BC0C96;
defparam prom_inst_5.INIT_RAM_20 = 256'hDC2FC6F09E70E71EF7234AE01EF3431BBAEF646E00046B3FFFEFFBFF9F4F1857;
defparam prom_inst_5.INIT_RAM_21 = 256'h8708FE60004D9DFFBEDFF887D98BFFFD8136FA15F7ADC3472D018A5D9AA5D4C4;
defparam prom_inst_5.INIT_RAM_22 = 256'h057BC75EFF39381813402A696B39E2E4D02A08BF0D5181F91DE87C93B9FA776E;
defparam prom_inst_5.INIT_RAM_23 = 256'h534C8DE6F4617B0CA1AB24FE2B14BB9B3B0E180C037A7FFDBFFE21E608FFFFB9;
defparam prom_inst_5.INIT_RAM_24 = 256'h2B0008005307FFE7FF85FDE8F03EEE0012EAD7B9A827B51E0F387492B0E2E725;
defparam prom_inst_5.INIT_RAM_25 = 256'h716AFB8060630700F6FA4CB774BABD8CA4F6E3ABB9FBDBCC15C01C1A9F1FF450;
defparam prom_inst_5.INIT_RAM_26 = 256'hF564C6C8399C51957200093077FC59AFC204083E595FFFFFFFFE0E134DF3E551;
defparam prom_inst_5.INIT_RAM_27 = 256'h040201F513FDFFF79FE7A1FDF8700FC79A8A6108233EAA4971A52AB8333FBAE4;
defparam prom_inst_5.INIT_RAM_28 = 256'hC41C0001F0B343C13318C645294AF2FBBA99671E077E132D000688D79F045A71;
defparam prom_inst_5.INIT_RAM_29 = 256'hCCCBC7F0F623B10001413FB7D1AD840010806EE12FFFF5E998082FEB2C2820FE;
defparam prom_inst_5.INIT_RAM_2A = 256'h0C1CDC5FFFA11C6633175F0EC1CD72244024000084EDE918CF8EC580AA945DA3;
defparam prom_inst_5.INIT_RAM_2B = 256'h4020035A88CEF9C7E3C849DC0CD9D9026CC5F23E34DABC072924FDF5725D0000;
defparam prom_inst_5.INIT_RAM_2C = 256'h617C076FA78F33147D996C541360000205C980FFFE68FF4468D1E3A0105E9108;
defparam prom_inst_5.INIT_RAM_2D = 256'h5B606FFFF8F6B541EE78F81022E8888144308B3497003D901FB12A0C7CA69B33;
defparam prom_inst_5.INIT_RAM_2E = 256'hFBD936592EA4009E069FFA8DB98B199C7C004E40F4F8EE3AD976293DBC000011;
defparam prom_inst_5.INIT_RAM_2F = 256'h001EC663E1D2EACEB3A9D84B0000845E6E1BFFBE3B6B7879EA1B2006EC400003;
defparam prom_inst_5.INIT_RAM_30 = 256'h84F9FFFA758283F78F080D9A0100457FD59F8A5A3B70327F0518C4EB919CCE7F;
defparam prom_inst_5.INIT_RAM_31 = 256'hC8E3CB0EF710FFBE38140B19D5771FD0036F132C8D2CBD5872BF31C002013C47;
defparam prom_inst_5.INIT_RAM_32 = 256'h43F95749DF6F6C0773172E45326E9E78FFFF7D7E0FD607E1D00030110005FDE1;
defparam prom_inst_5.INIT_RAM_33 = 256'hFFBE1F2DFE45F8DE20D051000057908646A9A0724F70639A6AE56BCF419FE046;
defparam prom_inst_5.INIT_RAM_34 = 256'hD8DEB35620BE05246BCA8671E7E0178BC4ABA78668DC63936E34C0407BF1980F;
defparam prom_inst_5.INIT_RAM_35 = 256'h751CC4D1761C64E6B71E026EFB5706FFF87F119D95FD3E80F3E000017260E458;
defparam prom_inst_5.INIT_RAM_36 = 256'hFE438EE9BF0FD8068009512FE02AC562F2F7F539F2F8D8B9488C7873E616FBF8;
defparam prom_inst_5.INIT_RAM_37 = 256'h44A558E88E0DA99E1ABC78F9820EA8488FDC97325D2059702D009BE59D81FF9F;
defparam prom_inst_5.INIT_RAM_38 = 256'hB1F9EB1FF1A2A2658FFFDCC1301FFF1FBD690BFFE5CF030D881457FC7B26C57F;
defparam prom_inst_5.INIT_RAM_39 = 256'h0C433F30E8802010080BC0CC7626D0048B14E882030F67F91C3C78806F44657A;
defparam prom_inst_5.INIT_RAM_3A = 256'hD7602D4A052901B05C2E0027E4DE6D8FFB333FF03780E865B4FC448C5FFFFFE7;
defparam prom_inst_5.INIT_RAM_3B = 256'hC20FFBED77282CFB7F322113FFFFFFC110CFFE2D0010001016FE2E120CF81E71;
defparam prom_inst_5.INIT_RAM_3C = 256'h0AFF8D4118000225FFCB8449580442129AFF18230896207C2F8067FF6B1BF14F;
defparam prom_inst_5.INIT_RAM_3D = 256'hF5041F827C07FA16441F7F708D995E270FFFF12845CF2329CF94A1FFFFE18E50;
defparam prom_inst_5.INIT_RAM_3E = 256'hFF8AB65D3B85F9B79D33FFBBF0BE4100D7E9A004100001DBA1C23FA93C1716EE;
defparam prom_inst_5.INIT_RAM_3F = 256'hFCC6A041790657D1F1A3F6C43678C72817F1800FBEF805E0191FFF873EF32707;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b1;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'hFC00C03CE307E007A7FFF0C7883A0FFFBACC3019D2F041614C3FEFFDBE28401F;
defparam prom_inst_6.INIT_RAM_01 = 256'hF9A416E3892998F303FFBE7C67EC2FFE3D802060000DD60E6E25602351A9383F;
defparam prom_inst_6.INIT_RAM_02 = 256'h07000120EFFFD6B954FFD1A4FE0C5B881CAE03000FB101FF7FFF80FD9583FDE7;
defparam prom_inst_6.INIT_RAM_03 = 256'h174C803BFE01E7EDF66F02AEC3FFB8FF956F0D61067628E06EF5FCE5C3866F9C;
defparam prom_inst_6.INIT_RAM_04 = 256'h61B41BBDFE7361FE7CFBA024DEDF24004400023BBF972644B0C416840C5F8201;
defparam prom_inst_6.INIT_RAM_05 = 256'h0C0016EFD9B9D577953F99D3BBE039FFFC0FFFBC1197DFFE8CFF83C26FFFCEC6;
defparam prom_inst_6.INIT_RAM_06 = 256'hDFFFB1000AFFFDF7EBFFF007FFBBE0D9C46DB7F873F43FFFFFE7C47BE1F8A800;
defparam prom_inst_6.INIT_RAM_07 = 256'h59636C0BC80FF9FFF1F0FFF47A3F6000000607F78A22BC8EBF0FEB07629DDFFF;
defparam prom_inst_6.INIT_RAM_08 = 256'h0401DEE3E6BDF45CF52D07D01FEFFFFFFF3C8004DEFF3DFA000001FFFEFF9CAA;
defparam prom_inst_6.INIT_RAM_09 = 256'hC200479FFFFAF800031203F7FFDB3EAA7980127B79BF9DFFCE6302FDCED00400;
defparam prom_inst_6.INIT_RAM_0A = 256'h058EAB723F7FFF1F88487FE1752015418E7FE038DB2DF00A9ACCF40FEEFFFFEF;
defparam prom_inst_6.INIT_RAM_0B = 256'hA1558B2D4204FBB8B6CC2F7A3F7FFF6080815BFFF77C0000029ECFB9FE3F36F5;
defparam prom_inst_6.INIT_RAM_0C = 256'h0036FFFDDF840001A68BEFFF8790915BA377ED4FFFFFDFFA140CF3FF0002308A;
defparam prom_inst_6.INIT_RAM_0D = 256'h6ED031F9B7FFFBE075FC3FC0000043BFFFE0F3274977E98407CF600FFFFFD810;
defparam prom_inst_6.INIT_RAM_0E = 256'h720A2D34EEE9981823E07C3CFC6000451BFFFDF3C07EE7E6B45FFFE078D6CCC7;
defparam prom_inst_6.INIT_RAM_0F = 256'h7FFF7CF82F7AD60676FBFF83C205FAD2F17A6DEBDC7EF8267FA5EC9023401C7F;
defparam prom_inst_6.INIT_RAM_10 = 256'h715FFE71FFFF285F30F85C82C04B1FBC80C4935F8DCC21CCE0D2033008014141;
defparam prom_inst_6.INIT_RAM_11 = 256'h0F1D0766C04CD93810081F0000007C7F9FFFFFFFFE3CA9ABFFFBF83F0ED2C826;
defparam prom_inst_6.INIT_RAM_12 = 256'hFFF5FEF0321F8CBFFFFF01BE64E9B0D947FBFFFFA72BFFF8FE00005E077FFF38;
defparam prom_inst_6.INIT_RAM_13 = 256'hBEEFFFE9E607FE3FC1002CA9C7EFBC80F1C70CC4FFA84D1000FC9000051F1FFF;
defparam prom_inst_6.INIT_RAM_14 = 256'h8E00C309959342083F23000007BE7FFFFFFEC94AD783AFFFFDDC01EC043FC672;
defparam prom_inst_6.INIT_RAM_15 = 256'h804CA86CCA1FFFFFFEC00C3880847E4F9E9F669EF3FFCFE022234A71FDEFFF07;
defparam prom_inst_6.INIT_RAM_16 = 256'hFFE7663C9FE36880007EF9FB9EFDC0585E93B8DAC4F80053EFA30000407DE7FF;
defparam prom_inst_6.INIT_RAM_17 = 256'h7C53771938000E103280C00E0FE840C301CFCFFC073FBFDE3F904839E393D3F9;
defparam prom_inst_6.INIT_RAM_18 = 256'hC038C3002FEFF7FDFD0E1A80E03B7BFFFFFBAE1BFA37A40135D9F8FA7FFB27E0;
defparam prom_inst_6.INIT_RAM_19 = 256'hFEF6D7FE3FDC10031BF7B7AFDFC81E0B4531320F800F8C3BB000001800399527;
defparam prom_inst_6.INIT_RAM_1A = 256'h049111E102A808030000009631523D79FC000019A6FFFDFBC842368DEA1FEFFF;
defparam prom_inst_6.INIT_RAM_1B = 256'hC000060807FF7EFE0A23FA7C8D7BFFF5D9A6FB8FE111072CFF77EBABDEC0E1C0;
defparam prom_inst_6.INIT_RAM_1C = 256'hFEDF83FE04C1D365D45ADB1FF43048F307E47880F203F9E00000321B2BFEC5F7;
defparam prom_inst_6.INIT_RAM_1D = 256'hCD1E003801C40C80013B7CA07FFFFECC000060008FFFFE03C06D91C75EFFFFFF;
defparam prom_inst_6.INIT_RAM_1E = 256'h0006FC2BFFFFFF1163E543EBFFFFFCD97DF0BFE11C266FEEA0FD9DD8C754BBB4;
defparam prom_inst_6.INIT_RAM_1F = 256'h7E5FE4C10183FF602BBD7FE0C5476B708F200F45F3810001187CE1FFEFFFFBC0;
defparam prom_inst_6.INIT_RAM_20 = 256'hC802D1FFE243F7F310D07FF8FF0107FEFE87C23FFFFFE66873116EFFFFFEB64B;
defparam prom_inst_6.INIT_RAM_21 = 256'hB173D3FFFFDEC8824397D7FE7FDFFFFF83F630A4016F900A2EFFCC27BB2A63A3;
defparam prom_inst_6.INIT_RAM_22 = 256'h6DAD1947D0777E13EFFC0CA08897087A00724FED0C07FBC8C00001235A6600ED;
defparam prom_inst_6.INIT_RAM_23 = 256'hE807FF93FE8844900004549FB70623126CE3FFFFF6C2E310C187BFDFFB7BCFC0;
defparam prom_inst_6.INIT_RAM_24 = 256'h12FFFFFFF9C45B276D7FFBFBFECFF83994620E0300E006F3BF83764DDE567E03;
defparam prom_inst_6.INIT_RAM_25 = 256'h10DC05805E03B0FFFC953C6BB70FE0D003FFC4FF728845000ECB7F7186AF8ECD;
defparam prom_inst_6.INIT_RAM_26 = 256'hEFD27CA31897803ADCEC6C79716765FBFFFFFFFFB86CA09B87B6FF7FBF70379F;
defparam prom_inst_6.INIT_RAM_27 = 256'hFFFDFEF2CF0859DFEFFFF790DF056C0051C3CCF11883EFFC662EAB1AC3CB4E40;
defparam prom_inst_6.INIT_RAM_28 = 256'hF082C3C4A3BFFF7AD22FC567733590377A3E3FBAC3E87BE80F30A21895A5D01F;
defparam prom_inst_6.INIT_RAM_29 = 256'hBF1C6B64A6F79333C037DF7945F0C56FFFCFFC5EE6E614CFFF7F3BBF80DBC05D;
defparam prom_inst_6.INIT_RAM_2A = 256'hFFFF43A44FC4639FFDEE7FC8EE8C064A81DA320C933F05D1F99610FFC8BF07F9;
defparam prom_inst_6.INIT_RAM_2B = 256'hC2E18204FBA35ECD6F0CBEE00DE2FF8E844BE06ECE255C0137E08C3358F92DD7;
defparam prom_inst_6.INIT_RAM_2C = 256'h0BF81FC82C74005DF70D7167551F7DCFFFF96334C7B027FD7BD4F10FDD110828;
defparam prom_inst_6.INIT_RAM_2D = 256'hFF356993D7E6BFFEE7FF07F84001FBBE80048337E3AB733EA42FD85B307FB801;
defparam prom_inst_6.INIT_RAM_2E = 256'h08604FE868630DD70FFEB96A0F1867ABFFFF158BF0007FFD1F0AAB2DB8717DFF;
defparam prom_inst_6.INIT_RAM_2F = 256'hFF189AE8001FFEA03AFC83C61DDDFFFF006D7FA5C8777FEFFF81CD400060A780;
defparam prom_inst_6.INIT_RAM_30 = 256'h15C0DA5D1FFF5DFFE00ECC417BBC98200011FC2C1B9AFBCBFF49BE578837A97F;
defparam prom_inst_6.INIT_RAM_31 = 256'h33FF03B4407480FD99BB93985F25FBFF2EE47800BFFC523B400037B90BFFFFF0;
defparam prom_inst_6.INIT_RAM_32 = 256'h95600007BE11BB000060A72FBFFFE89CBEE06F80BFF60E7C0FF0022E2E841000;
defparam prom_inst_6.INIT_RAM_33 = 256'h000E6C2FFF92DF28F0004BAB01E0200DB60C2DEC6240FFF00FE45E5AF67FFF2D;
defparam prom_inst_6.INIT_RAM_34 = 256'h42653DA371BFFE27F6547FBA5FFF7CF0E63901CF3023C000198411AFFFFBE9AF;
defparam prom_inst_6.INIT_RAM_35 = 256'h88000C0A2070200060C08577FFEC7BA55C9AC767BF77A2BF7012E080671003FE;
defparam prom_inst_6.INIT_RAM_36 = 256'h9090FFF9DFE01FD100246006800035D9B850329C3FFFF17EF415951F7F730FF9;
defparam prom_inst_6.INIT_RAM_37 = 256'hB5F98F3FFFFBFFFF8CB78FFE7C89FE4000010466B88000078E1FE7FAFC05BD2C;
defparam prom_inst_6.INIT_RAM_38 = 256'h0003705E800007E0C529FDB3400B7789C539FFFFF00FED955B10566208F7EBD4;
defparam prom_inst_6.INIT_RAM_39 = 256'h667FFFFC017DE454C19D18820FF4EF2E4C8783FFFFFFFFE4BCC7FE5711FF8800;
defparam prom_inst_6.INIT_RAM_3A = 256'hD1811FFDB7FFC28E67FF55F27FE04100004A5E000000F036C7B3F280183DD2D9;
defparam prom_inst_6.INIT_RAM_3B = 256'h143F800000202158FFFF0802066D50577F7FF628FF234001A2E786FFFE756F7E;
defparam prom_inst_6.INIT_RAM_3C = 256'h3FFCC21F1D85E3BDB1FA1FFA1B2856127037FFFFED99B031F628F1FFF6000000;
defparam prom_inst_6.INIT_RAM_3D = 256'h03FFBFFFE98FD87F1141FFFFA000003A90FC2000200027A7BCC000830130759C;
defparam prom_inst_6.INIT_RAM_3E = 256'hDFE00000801FE904C0003ABC1BFEB07BA7F107F3008666EF6203DE8180D47530;
defparam prom_inst_6.INIT_RAM_3F = 256'hFC40FF969DF8F3B73FFFE2773DAD1E07EFFFFFF0DE881CB520FFFBE0008006C0;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b1;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'hFFFFFC68E6071FE7BFFFF84110011CDFF871382807255100010F1F90DDBA1EF5;
defparam prom_inst_7.INIT_RAM_01 = 256'h04800000D5D9918003DEB556ACC03F9F86FFD6AEEFF9F9DBFBC3EA8BF1A787FD;
defparam prom_inst_7.INIT_RAM_02 = 256'h03F96FB757FFFFFF0194EE1B91C073FFFFF41565902DB9BFFFFF810001DFF3FE;
defparam prom_inst_7.INIT_RAM_03 = 256'hD0034FF109FC79FFFFFE100C32487F7D93000019AE203037EA9533178C06A840;
defparam prom_inst_7.INIT_RAM_04 = 256'h400007AC60000CFFC8F26309016F20C75F17EFFBFFFFFFF9931D347DC811E73D;
defparam prom_inst_7.INIT_RAM_05 = 256'h42FFFCFFFD9FEC491FB4927019F9AFF4055F600DC01FFFFFFFE4001C5ADFF684;
defparam prom_inst_7.INIT_RAM_06 = 256'h5D500F918043FFFF7B002F66E3FA7FF004015A7600002FF3EE8B0308423C03EA;
defparam prom_inst_7.INIT_RAM_07 = 256'h0266F7200037FEA0ECA67608A00E7EBFFFFEFFFFFFEE22DB0173D808C6D87C56;
defparam prom_inst_7.INIT_RAM_08 = 256'h7FFFFDFFB836E4F6D6C600A9D40F3BB9A803D0201081EFFFF87BE1F9FFFFFC47;
defparam prom_inst_7.INIT_RAM_09 = 256'h07A4F1015FE9E7F432DA0F5FFFF691921F2191000FEFDB440D55E01D030DF3BE;
defparam prom_inst_7.INIT_RAM_0A = 256'hC0D0010CFF27807CAD95604001FF6FFFFFFDFFF433D4F1AD73E0180219005306;
defparam prom_inst_7.INIT_RAM_0B = 256'hFFFF9812037E7F0DC180068000BF21A0F3060401F3FFFC043E5357FFFFEF9C5F;
defparam prom_inst_7.INIT_RAM_0C = 256'h5581001B7DFF010F9DF8FFFFE37F09F4A0F4833F9652F8682981003274EEE7FF;
defparam prom_inst_7.INIT_RAM_0D = 256'h7828FFEFD77075E118901C3FBACFFFFF9FFA0B77F9E67B10000380402454C7EF;
defparam prom_inst_7.INIT_RAM_0E = 256'hBF8927F5B782980018004432FA71761E8408007FFFBA26E7423FE7F5FFE1FC7A;
defparam prom_inst_7.INIT_RAM_0F = 256'h10501FFFFF83B06CC7FFD3FF6D1B0A2F254FEFDC83374A66C0256DCF3F87FFE9;
defparam prom_inst_7.INIT_RAM_10 = 256'h5EFFFF00D73D1450034277BFDFFB1FEA8159D78FB5050002000E4B2E9EDD1171;
defparam prom_inst_7.INIT_RAM_11 = 256'hB4AD399651C00000008345DFBF288D040007FFFBE3BF2E84FF8E9FBB7ECEA7C8;
defparam prom_inst_7.INIT_RAM_12 = 256'h221D7FFF39E181FEAFFBFDFEF5617CDEFFFF8A30ED2EEA00F06DFF6EBF5EFA8C;
defparam prom_inst_7.INIT_RAM_13 = 256'hFFB987EE84D5E04527E77FBFBFF0837B504C39E470000800066A937EA2561000;
defparam prom_inst_7.INIT_RAM_14 = 256'h94074D1C00000006FBE9EF4C65E4101C273FFFCEBDC4EDDDF8FF7FED2FAFFBFF;
defparam prom_inst_7.INIT_RAM_15 = 256'h81FFFB0F6BFA73FF98FFFA62C7FE3FFEEB14C4E96CEEBF32FCFFEFF8C038896D;
defparam prom_inst_7.INIT_RAM_16 = 256'h86C54188B7FBE0AFF77FFE0073EFD7CF18EA8E800000187654FFD95A78800080;
defparam prom_inst_7.INIT_RAM_17 = 256'hBCA3E200002019717FCC3D3FB014000817DEF7357F6E6CBFBF7FBD5FFFFFFFEF;
defparam prom_inst_7.INIT_RAM_18 = 256'hFFFECAC5FFFD2BEFC7CD18FFFFDFEBE0D144715C7FF01FFFFFFF80230FAC75FC;
defparam prom_inst_7.INIT_RAM_19 = 256'h8F5CAF1FFC17E6F7FFE0F602C48808A238FF00000206A05FF5E94FED04000201;
defparam prom_inst_7.INIT_RAM_1A = 256'h2C000402133197F8102786084101A03EEF0BD5A07C0A5E79F362B7FFFBF4383B;
defparam prom_inst_7.INIT_RAM_1B = 256'hF89A1DAD01F9C9F66E9FFBFFFED802379D26242701FFFFFFD87ABD05CFB8C0AB;
defparam prom_inst_7.INIT_RAM_1C = 256'h5C44B9E15BFF85543CE273E5845C8EE64000021E2C73FD688ADF91A0000900CF;
defparam prom_inst_7.INIT_RAM_1D = 256'h011001CF7DFFD136B7986100000003FC3BDFD7F87E77CA4E9B3FF7FFA600FFBD;
defparam prom_inst_7.INIT_RAM_1E = 256'hCDB9F1F0FFE2A315FFFF79600050CF1295EC182BFBFF7F1CA43BD1D516BD59B4;
defparam prom_inst_7.INIT_RAM_1F = 256'h5C040FFEBFFB0CBF0C79D51D80D779F9607354227E2D029D8601600182082BCF;
defparam prom_inst_7.INIT_RAM_20 = 256'h9FFBD27D1AD5A7FFE2340660820AF7F3C867818E48E6457CFA9948000EF043D9;
defparam prom_inst_7.INIT_RAM_21 = 256'h6A5DB3505E36A073FCC00812DD8EB3BE4A013FFFFF8F702329E0A3734AE6E639;
defparam prom_inst_7.INIT_RAM_22 = 256'h00B8FFDDDBBF5946A14C9D3CB1AFF19DFCB3DF2F8830FFD81F5F6C0E8007FCD3;
defparam prom_inst_7.INIT_RAM_23 = 256'h3CE306DCCCBFFE8FFFDFF8F0007078E39E5F01C57C428F294004187E721123AC;
defparam prom_inst_7.INIT_RAM_24 = 256'h9D2F6A5D3093090000C61F36D65DA40F0F7FEFC0D904782B9672DF047FFBFFFD;
defparam prom_inst_7.INIT_RAM_25 = 256'hDFFFF0B52C60417107E9651FF71FFB5488C17FF00FFDFBBFFFFFFFFFDFFFDD74;
defparam prom_inst_7.INIT_RAM_26 = 256'h00D259CBBBF17FFFF5DCFAF7258527A2968153140CD900014987E39BBAD3E3C3;
defparam prom_inst_7.INIT_RAM_27 = 256'hA5813EC3C004000413D393FAB9DE2237FB7C1A6A69A05695E620D3FFFFFFD6DC;
defparam prom_inst_7.INIT_RAM_28 = 256'hEF2D8614E0281EFF380817FF7DE4C13C70A6E2AFFFFF7E75E58908D20FE88BB6;
defparam prom_inst_7.INIT_RAM_29 = 256'h70B8BBFEFFFB6C002FBE0201463F5717AF1F80C04080110D3D658015EF673F7F;
defparam prom_inst_7.INIT_RAM_2A = 256'h932110001159E3FFD04046519C03D3E587E78B382E8CCDD43605FFDFF8FD8C72;
defparam prom_inst_7.INIT_RAM_2B = 256'hF4FE4A00F1F84E9183FF7F9825200862E0067FFFDD06A01D83C0FE5F54AFAE50;
defparam prom_inst_7.INIT_RAM_2C = 256'h80BEFC7B0001FCB19A9BBECAAD76081EA84A4008678F7FEBC83C7F6F803BD067;
defparam prom_inst_7.INIT_RAM_2D = 256'h0002013C2BFBDDBC8384A2C00BFC0844F2552B8D39639F697BFFFE02B40E441B;
defparam prom_inst_7.INIT_RAM_2E = 256'hFDA701D824139C1FFFFF80F4425B7E6801FDFE0200FEA59D8BFD844D9F1401FF;
defparam prom_inst_7.INIT_RAM_2F = 256'h78384025D4B236CA1ED28B183E2103E101CFFF765EFFF32C1FF2F81FB060D5EA;
defparam prom_inst_7.INIT_RAM_30 = 256'h33FFFAFFDFFC747BE03682A10813643D206CA78032130A7FFF25D91B8F9DAE40;
defparam prom_inst_7.INIT_RAM_31 = 256'h14132BD4E924E7FFCA9A8962A56B82160E10096C23766BAD1166A4AFD003FC90;
defparam prom_inst_7.INIT_RAM_32 = 256'h40BC78F77DA6CA08451D01F8127DC83F7FEFFFFFDD588132016827223B8C8E48;
defparam prom_inst_7.INIT_RAM_33 = 256'hEDDFFFBFF4673F86C00A003863B7BC40971618AAB087FE620DA2E9A353E10140;
defparam prom_inst_7.INIT_RAM_34 = 256'h875C3C9E01848C243B3C7B6CFC11002061FE326A0CA9E52ECBF85FC859A9D629;
defparam prom_inst_7.INIT_RAM_35 = 256'hEE39AB9C0E1EDB34D80FF21ADB9FDBAAFFF1F7FD4387E89E04805FDBC9CBE641;
defparam prom_inst_7.INIT_RAM_36 = 256'hF9FE776393C91B8240193F8284938706C75447062124825BFC115A3F00000009;
defparam prom_inst_7.INIT_RAM_37 = 256'hFEB7C0578803D7FF475817F00440007B0CD757976B71E8B6881D0397C77FCFC3;
defparam prom_inst_7.INIT_RAM_38 = 256'h78293E3497639F3012D825F3FFF3F5D67E7DDE9F7BC390503D5EB125449149A6;
defparam prom_inst_7.INIT_RAM_39 = 256'h3F95C9DB78F6743AF14AE10AFA66B96130705500285677D76EF1F400006147DA;
defparam prom_inst_7.INIT_RAM_3A = 256'h38408100327F19931CEE0000082F870123C71D68949D08027800CE7BFFEFE7FE;
defparam prom_inst_7.INIT_RAM_3B = 256'h051609B047F8B0FF1887FFFEA97E7606FEF072471FB85EB43CAA2385FFAC1C94;
defparam prom_inst_7.INIT_RAM_3C = 256'hFCC86B27E6FC048EA02E7D9EB314D03E1000027977FA6A8B1BC4001045E19A21;
defparam prom_inst_7.INIT_RAM_3D = 256'h00085F95B0D87AC2F0480471F4CD76423515217561063E6601FEFF38B433803F;
defparam prom_inst_7.INIT_RAM_3E = 256'hBC1D527B1D901C820FFFF7E3CAE6C74F143A12FA7C3DD372E58BABFC3EA2FF98;
defparam prom_inst_7.INIT_RAM_3F = 256'h0000F7BF015E1B207950DF4D7563FC000001443B068B10FDC0127FF9466729C7;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b1;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'h0000000931EDFFFFFFFFFFFFFFFFBFFFFFFF679FFFFFFFFFBFFB210000800BF7;
defparam prom_inst_8.INIT_RAM_01 = 256'hBFFFFFFFFFFFFFEFA15007840004FFDBFE54600000C00000037FEFFFFB800000;
defparam prom_inst_8.INIT_RAM_02 = 256'h97C0C80328020000DFFFFFF600000000000000403F7EFFFF767FFDFF87DBFFFF;
defparam prom_inst_8.INIT_RAM_03 = 256'h000021597FFFFFFFFFFFFCFFBA7FFFFFDC6DBFFFFFFFFFFFF9500040003FCFED;
defparam prom_inst_8.INIT_RAM_04 = 256'hE7DDD7FFFFFFFFFFF45960000177F7E4C06E020000000077FFFFFE1000004800;
defparam prom_inst_8.INIT_RAM_05 = 256'h80013000000C3F7FFFFEC00000678000000001397DFFF9FFFFFFC819F61D8007;
defparam prom_inst_8.INIT_RAM_06 = 256'h0000184EF7FE79FFFF300210006001999A76FFFFFFFFFFFE8E22000076FFBA01;
defparam prom_inst_8.INIT_RAM_07 = 256'hE0FCFFFFFFFFFEDFFA084003FFFC80000044000003FFFFFFFED0000021880000;
defparam prom_inst_8.INIT_RAM_08 = 256'h00000022DFFFFFBE4000002E1060000000021B79DFFFFF4C0208100108032B43;
defparam prom_inst_8.INIT_RAM_09 = 256'h0100637FB41E8600000040400B664A2D02CFFFFFFFFFFFFF0610007FDB020002;
defparam prom_inst_8.INIT_RAM_0A = 256'hBFFFFFFFFFFFFFF992001FF700001000000020F3FFFFB2080000544800000000;
defparam prom_inst_8.INIT_RAM_0B = 256'h20063CFFFFEF420000183515C00000005818FFE807A0800008205002C86A8860;
defparam prom_inst_8.INIT_RAM_0C = 256'h01FF8696003008200000001049C0027FFFFFFFFFFFF7FAA10003F8C100000000;
defparam prom_inst_8.INIT_RAM_0D = 256'hFFFFFFF7FFFFACD400DFC4000000000018B3FFFFFF7400000B07212B00000000;
defparam prom_inst_8.INIT_RAM_0E = 256'h27FFFFFFFB0000033BD0C3E0000108007FE020800C0100000000001A800037FF;
defparam prom_inst_8.INIT_RAM_0F = 256'hFE068000000200000000184E081FFFFFFFFFFFFFFFE3F4300F50444000000010;
defparam prom_inst_8.INIT_RAM_10 = 256'hFFFFFFFFF593C817C02000000000011DEFFFFEF340000CA70B3200000000241F;
defparam prom_inst_8.INIT_RAM_11 = 256'hFFFFFD008007F989E7003000100539F786440C000000002000038AEF0DFCFFFF;
defparam prom_inst_8.INIT_RAM_12 = 256'h910300000000000000622DC1FFFFFFFFFFFFFFFD7CFC0060000000000002803F;
defparam prom_inst_8.INIT_RAM_13 = 256'hFFFFFFF7FB8030000000000001003FFFFFBB40400804039E8010A04100CFFBE1;
defparam prom_inst_8.INIT_RAM_14 = 256'hFFA4000C0007E380238007F9FE7FDB837000000000001080009D1C73FFFFFFFF;
defparam prom_inst_8.INIT_RAM_15 = 256'h10000C000008000001844F5FFFFFFFFFFEFFFB87FA0BC10000000000200FFFFF;
defparam prom_inst_8.INIT_RAM_16 = 256'hFBFFFEFFC2048000000000141FFFFFFFFE000E001236C0E0693FF7DFFFFDF962;
defparam prom_inst_8.INIT_RAM_17 = 256'h80020912EEBC326E5FFFFFFFFEEFF88000F000000000000042EC5FEFFFEFEFFF;
defparam prom_inst_8.INIT_RAM_18 = 256'h0240018100000000F8FFFDFFFFEFFFFFFFFFFFF08000400000000D877FFFFFEF;
defparam prom_inst_8.INIT_RAM_19 = 256'hFFFFFF00000010000002877BFFFFFB68040001C14B005840FFFFFFEFFF7A0000;
defparam prom_inst_8.INIT_RAM_1A = 256'h1200637ADE1D640FFFEFFFFFE6C00000000068400000602233FFFFBFFFBFFFFF;
defparam prom_inst_8.INIT_RAM_1B = 256'h0000800000003D3FDAFFFFFFFFFFFFFFF77FC0000004000000D0EEFFFFFEC400;
defparam prom_inst_8.INIT_RAM_1C = 256'hFFB400000000000001FFFFFFFBF1261141613465B95C02FDFFFFFFFE60000000;
defparam prom_inst_8.INIT_RAM_1D = 256'h3D4F8ADFAD807BFFFFFFFFE00000000101010000000B0EFFCFFFFFFF7FFFFFFF;
defparam prom_inst_8.INIT_RAM_1E = 256'hC0A0000002C3FFDFDFEFFFDFFFFFFFFFFE02000000000000A7FFFFFFEB60959C;
defparam prom_inst_8.INIT_RAM_1F = 256'hC040000000000045FFFFFFFBF180717833F92C0B2401FFFFFFFFF8000000FF01;
defparam prom_inst_8.INIT_RAM_20 = 256'h7D76B77F5B5FFFFFFF7618000BF761400055002020FFAFFFF7FFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_21 = 256'h0100004F97DFFFFFFFFF7FFFFFFFEFD01000000000008DDFFFFFEFFC000618FF;
defparam prom_inst_8.INIT_RAM_22 = 256'h040000000000EFFFFFFFBF8800E93FDFF54C8FF23FFFFFFFF4800005FB3C8200;
defparam prom_inst_8.INIT_RAM_23 = 256'h2E4FCB3CFFFFFFF6400001E5C51C000025010307FBFFFBFFFFFFFFFFFFFF7C00;
defparam prom_inst_8.INIT_RAM_24 = 256'h40016FDFDBFFFFFFFBFFFFFFFFFF808000000000201F6FFFFFFBE00008A7FFED;
defparam prom_inst_8.INIT_RAM_25 = 256'h00000068FD79FFFFF3C8025F097FFEB3C1DF13FFFFFFFF4000039F0EA5800000;
defparam prom_inst_8.INIT_RAM_26 = 256'h5F86E367FFFE480003800447600000100269F7F9FBFDFFEFFFF7FFFFFFC00000;
defparam prom_inst_8.INIT_RAM_27 = 256'h000FFDFFF77B3FE7FFFFFFFFF00000000000045FFFFFFFFCD20000C937F61BF2;
defparam prom_inst_8.INIT_RAM_28 = 256'h00007FFCFFFF3FE9E02FFA62FEC2FDA66BF7FFFFFFF000204424C7D600000400;
defparam prom_inst_8.INIT_RAM_29 = 256'h0D48BFFFFC80003845362360000000000EDFFFBCFCD97FFFFFFFFFFC20000000;
defparam prom_inst_8.INIT_RAM_2A = 256'h87FFFF3F33DFFFFDFFFFFF00000000040001DFFFFFFFFFD90275FFB1A2FFFB84;
defparam prom_inst_8.INIT_RAM_2B = 256'h006BFBFFFFFF0006AE7FBC77FFFF7D07001EFFFD20001B9DAE823E0000000003;
defparam prom_inst_8.INIT_RAM_2C = 256'h01DFFFA0000653E80CC590000000001EEFFE7FF7B9FFFBFFFFFFC00000000001;
defparam prom_inst_8.INIT_RAM_2D = 256'hF3FFFFBFEEDFFFFFFFF00400000002316F7FFFFFFFEBC7234FFC94FFFFEEA060;
defparam prom_inst_8.INIT_RAM_2E = 256'hFFBFFFFFFD9A70FFFF068FFFFAD05C002B7FD60043C46179C83C00000000003C;
defparam prom_inst_8.INIT_RAM_2F = 256'hFFE60200F8EDBF76F700000000000C3E7FDBDDFBF1FFFFFFFC00000000000677;
defparam prom_inst_8.INIT_RAM_30 = 256'hB7FEFFEEFFFDFFFF00000000000917FFFFFFFFFFF8F3BFFF983BFFFF58478001;
defparam prom_inst_8.INIT_RAM_31 = 256'h7FFFFFFA005B7FC6263FF9E741A00005FD40003E96BFEEF6F00000000000BF3F;
defparam prom_inst_8.INIT_RAM_32 = 256'hD0203FD3DFFBA61D00005880001FCFFFE6BEFBDFFFFFFFC0000000010D8BDFFF;
defparam prom_inst_8.INIT_RAM_33 = 256'h9EFE7FFFF7FFF00000000043E6B77BFFFFFFF7A11F7FF9874BFF43E1DE0001FF;
defparam prom_inst_8.INIT_RAM_34 = 256'hFFFF61F8FFD70E273C68E083FA003FF800017A9FF5B84F80001DEA01004DFFFB;
defparam prom_inst_8.INIT_RAM_35 = 256'h00163E483846780008001080C3EEF597FCFFFEFFFBFC00000000042FFE5FFFFF;
defparam prom_inst_8.INIT_RAM_36 = 256'h6167FDFFFF0000000010127BFFFFBFFFFFFCDFCFF4BFF347D48C4EFF801FFFC0;
defparam prom_inst_8.INIT_RAM_37 = 256'hFE29DAF85FFE1C2E2ACB5FF807FFF00047D2576F9C3E000580062433F8BFE3FE;
defparam prom_inst_8.INIT_RAM_38 = 256'hF22B45D02FA00026020026DCFDFBF7FCDF7FFBFFC080000004055EFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_39 = 256'hFFFEFFF00000080013FFFF7FFFFFFFFD7281A35BFFFCFF0194A07F01FDDC284F;
defparam prom_inst_8.INIT_RAM_3A = 256'h48A37FDFFE6F20F7500FE0FFFF5D73FE6D902101780000002001A37FFF4FFFAF;
defparam prom_inst_8.INIT_RAM_3B = 256'h8740A0BF000000002037FFEFE77FA7E76B3FFC00000000007BA767FFFFFFFE45;
defparam prom_inst_8.INIT_RAM_3C = 256'hFDFF000000011201DFFFFFFFFFFFCAB20413FFBF92800A9780F83FFFFFDDFF82;
defparam prom_inst_8.INIT_RAM_3D = 256'h1B0FFFEB8003877B3F03FFFFFFFFF93FF04345F00000000058CCFFFE19E76E1B;
defparam prom_inst_8.INIT_RAM_3E = 256'h2B81FC0000000026333FFF9E79D9E3FF7FC000000005287BCFFFFFFFFFA646C0;
defparam prom_inst_8.INIT_RAM_3F = 256'hF080000204D21F6EDFFFFFFFECFA1819DFFFDFAC4473E70F807FFFFFFFFEA8FA;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b1;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'h3FFF8F0541F4F0C03FFFE81A3FE2C343024BC00000800B40FEF5F87E4423314F;
defparam prom_inst_9.INIT_RAM_01 = 256'hC9700000000037FEFFBFE7E3F93D77FC000000103ACEFD7FFFFFFFD83AE901CE;
defparam prom_inst_9.INIT_RAM_02 = 256'h00004916463707BFFFFFFC836B900F6BC5A903EADE3E3803FFE7275F3E62E90E;
defparam prom_inst_9.INIT_RAM_03 = 256'h4080B70EC39C00FE023CFA53CC9E0CE03F0000000004FF9FEB79F167BEFF6F00;
defparam prom_inst_9.INIT_RAM_04 = 256'hE0000000848EBDFFFFF03877DFDFC0000000011187B2CFFFFFFF217750161436;
defparam prom_inst_9.INIT_RAM_05 = 256'h0009023ADC3871FFFE0010F829D90D6027CB4748E7400E08CA8C0C0082EC57FF;
defparam prom_inst_9.INIT_RAM_06 = 256'hDB17C33BC0000CA8665030712D2E68FE00000002236F779F7B873FF9FFF04000;
defparam prom_inst_9.INIT_RAM_07 = 256'h000000015FFFDEFE40817EFFFC000000030002010361FFFE80141D31FB1C1C0F;
defparam prom_inst_9.INIT_RAM_08 = 256'h601B898428FFF4B401816329B7F003FA25BF44F00005017FDA6FB220F56D87E0;
defparam prom_inst_9.INIT_RAM_09 = 256'hCCD2380025AA62A99244D533FF9EFC000000003FFDFFFFF967FFFFFF00000004;
defparam prom_inst_9.INIT_RAM_0A = 256'h000C3FFFFFFFE6187FFFFFC00000002401000001E17FFE03A050A887E400348F;
defparam prom_inst_9.INIT_RAM_0B = 256'h680000B09EFF01EA1652EDFF00161EEE349F800E8B1B7CD6D6CB53E79BEF8000;
defparam prom_inst_9.INIT_RAM_0C = 256'h47A007751FFCAC0A5B4ACFCFF2F02000002DFFFFF8E011F978DEF80000000019;
defparam prom_inst_9.INIT_RAM_0D = 256'h13FFDF9E7F1AED1FFF7E00000000810100311382B08074A5068BFF003A0DAC6D;
defparam prom_inst_9.INIT_RAM_0E = 256'h5B6064B04C1CDA00817EF80D5776B3A3E803B04613CF3D3F2ECB2D8BBF400100;
defparam prom_inst_9.INIT_RAM_0F = 256'h01D2AD2FF9863B15D3170731F00000009FF7FFDF9F78A7EFFF20000000000400;
defparam prom_inst_9.INIT_RAM_10 = 256'hDFFFFDE7A0F8DDFFC00000100000200CAA0F9C820795301A878C0095E35C78FC;
defparam prom_inst_9.INIT_RAM_11 = 256'h80382B81DC7D008AF1CA34BA3F787E80F96A8781EAEFD7FC5E79F7BFFB0003DF;
defparam prom_inst_9.INIT_RAM_12 = 256'h8B8380066CA577AC7E0981FE4200FFF4FFFEFFF90F375FF00000000000000A71;
defparam prom_inst_9.INIT_RAM_13 = 256'hFFFFF3847F7DFC00100008100002FF60EB1FE0761E002D8046D2D73FBE3FA03A;
defparam prom_inst_9.INIT_RAM_14 = 256'hF6D01E006B03364172BDFFDE6BF01D45E383F06BFC46FC5E3BDFC7D023CFDEFE;
defparam prom_inst_9.INIT_RAM_15 = 256'hC3FF86C6B9C7AF0451E03ECCF3F7FFFFFFE69118FEFF000000000000C860B6D2;
defparam prom_inst_9.INIT_RAM_16 = 256'hF932481FFFC8000000000019A1240550461F9CF38BC18D945CDE3E48FC066BD4;
defparam prom_inst_9.INIT_RAM_17 = 256'h05F21C2289589162AF81FB3F07E5C740FFF85B827C35A35EB403B33EFFFEDFF3;
defparam prom_inst_9.INIT_RAM_18 = 256'hFF8BA79F41F5AE5E00D3FFFF35F9FCFEEFBCEFFFF000000000000E102302B077;
defparam prom_inst_9.INIT_RAM_19 = 256'h707BFFFD800000000007761580492043E067C1F414540EB3DC3CC3E7EB37D07F;
defparam prom_inst_9.INIT_RAM_1A = 256'h5D6C3B922C03E7FBF939FBFB78CE37FFF97BFF72159FD5AFE2BFFCFBFBFFF859;
defparam prom_inst_9.INIT_RAM_1B = 256'h2F56C60E8F790FFCF9FFFEF7FFDE7E603FEFFFB400000040017F020F41EB41E0;
defparam prom_inst_9.INIT_RAM_1C = 256'hFBDFF000000000005D77A2409A30F1E9FC81203381FFFF0ECE7FFCE2DB0FFFFF;
defparam prom_inst_9.INIT_RAM_1D = 256'hD88600084CFEF7330FFFBADCC1FFFFC89CD0C98228E301F27FBEDFF7E1FBBA82;
defparam prom_inst_9.INIT_RAM_1E = 256'h221D128C82000D47FFBBFC99DE975030F7F0000000000217B734756B0C38740F;
defparam prom_inst_9.INIT_RAM_1F = 256'hFEE00000000000006812FE3A3E7368E61084C010BF3A1987FFEA68B0FFFFF157;
defparam prom_inst_9.INIT_RAM_20 = 256'h200C36DF800C60FEFA7A261FFFFC731A82EB426E0004E5FFFFEFFBFF9F4F1877;
defparam prom_inst_9.INIT_RAM_21 = 256'hD8FC3E00005CCFFFBEDFF887D98BFFFF8100000000000174400FF65E1CC9DEC2;
defparam prom_inst_9.INIT_RAM_22 = 256'h00000000000033E01FBFBB8E723B2056075DE34F03307FFE61A503FFFE344C20;
defparam prom_inst_9.INIT_RAM_23 = 256'h6C72C661CC1FFBDA5164FFFFCE210810290E000003E9FFFDBFFE21E608FFFFF9;
defparam prom_inst_9.INIT_RAM_24 = 256'h730008007F7FFFE7FF85FDE8F03FFE00000000000007C81DF0FB871CC02215F8;
defparam prom_inst_9.INIT_RAM_25 = 256'h01000000404C07F877038F380DC401135AA110E787FBE0A86C3FFFE25FC206E0;
defparam prom_inst_9.INIT_RAM_26 = 256'h8D9C21C7F99EF0BF0DFFF1FEEC80BD17C000083ED7FFFFFFFFFE0E134DFFE400;
defparam prom_inst_9.INIT_RAM_27 = 256'h000201D0FFFDFFF79FE7A1FDFF7000000000000825E30C012D47CB47F410249B;
defparam prom_inst_9.INIT_RAM_28 = 256'h0000000045F03F38C3E0F9FF30460D20C678E0FE07A35762FFF8CD4AC02D8EF0;
defparam prom_inst_9.INIT_RAM_29 = 256'hBC383FF0E787C8FFFE6BFD901BCACC000080629FFFFFF5E998082FFFEC200000;
defparam prom_inst_9.INIT_RAM_2A = 256'h0C16C3FFFFA11C6633075FFEC00000000004000183A4F720F00FC7B1104BA43F;
defparam prom_inst_9.INIT_RAM_2B = 256'h40200311E2BC51F803C069801F241F1E1C3FF238F95D83F83855CC06E4F70000;
defparam prom_inst_9.INIT_RAM_2C = 256'h1FFC07A38CE0CC61BEFC10BBBC60000207987FFFFE68FF4468D1FFA020000000;
defparam prom_inst_9.INIT_RAM_2D = 256'hCB1FFFFFF8F6B541EE7FF810000000014430FC61A387C000000080070206870F;
defparam prom_inst_9.INIT_RAM_2E = 256'hFBEE394933040001F973E0B219870783FC0077388C004C6B670938FADC000011;
defparam prom_inst_9.INIT_RAM_2F = 256'h001C216DE1A1E25F8C0C6AC300008479E1FFFFBE3B6B7879FFFB200000000003;
defparam prom_inst_9.INIT_RAM_30 = 256'h7FF9FFFA758281F7FF0804000100457FF8EDF460DFF00FFFFDD86BCF8F83C1FF;
defparam prom_inst_9.INIT_RAM_31 = 256'hBE6E8D0C0B0FFFBFDA899C87C3F0FFD003A9A1D33E3373C7836488E000013C30;
defparam prom_inst_9.INIT_RAM_32 = 256'h76A492F6E35CA3F851D60E00027EC607FFFF7D7E07D637FFD00000100005FFFE;
defparam prom_inst_9.INIT_RAM_33 = 256'hFFBE1F2DFE45FFFE200041000057FF5B1BF656F1C3F003F393DEE7C0C07FE000;
defparam prom_inst_9.INIT_RAM_34 = 256'hD4ECCF31E000063A39C781F01FE0000D29DFF40440F3FC181554C0007F8E87FF;
defparam prom_inst_9.INIT_RAM_35 = 256'h1E15EED191FF867C9B3A027FE1B0FFFFF87F119D97FFFE800000000173FF06CF;
defparam prom_inst_9.INIT_RAM_36 = 256'hFE438EE9BFFFD8000009512FFFC138E906B06CF80C00E0D58783F80FE60003A8;
defparam prom_inst_9.INIT_RAM_37 = 256'hBD933817700FEEDE05FC07F98000B482C062EA51FFF8A4466880FFCD047FFF9F;
defparam prom_inst_9.INIT_RAM_38 = 256'h788E58FFFE3628BC4FFFC5BB0FFFFF1FBD690BFFF9CB0004081457FF82322900;
defparam prom_inst_9.INIT_RAM_39 = 256'h0C423F3FF8800000000BFF30665C2FD9B68C17FDFC054806FC03F8800006F45F;
defparam prom_inst_9.INIT_RAM_3A = 256'hB31FFFFFFCF1FFF003FE000000F5ED25E790FFFFC54DB3221482DE43FFFFFFE7;
defparam prom_inst_9.INIT_RAM_3B = 256'hA1FFFBF1AFB55584839890FFFFFFFFC110CFFFFD0000000016FFD01E868FFC54;
defparam prom_inst_9.INIT_RAM_3C = 256'h0AFFFF4110000225FF740677A7FDB74987FF1820FF162003FF8000000CBDC1D0;
defparam prom_inst_9.INIT_RAM_3D = 256'hF504007F800005FFC4000000EB738760FFFFFE35E5BAD173356C5FFFFFE18E50;
defparam prom_inst_9.INIT_RAM_3E = 256'hFF8B44FD7546818C470DFFBBF0BE4100D7FFA000000001DFFE03860EC79A5261;
defparam prom_inst_9.INIT_RAM_3F = 256'hFFC6A000010657FE01CFE068D4D5A0E8000E7FF00007FFE00000000640EE60FF;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b1;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'h03FFFFC31CFFE000000000F80F99FFFFBAF0E4657F5C402DC3FFEFFDBE28401F;
defparam prom_inst_10.INIT_RAM_01 = 256'hFE3EA17A0FA387F0FFFFBE7C67EC2FFFFD800040000FFFF0738CB8D75B18F800;
defparam prom_inst_10.INIT_RAM_02 = 256'h07000100EFFFE83E6390F8DAA67C0477FFFFFEFFFFB00000000000FE0C7FFDE7;
defparam prom_inst_10.INIT_RAM_03 = 256'hFFFF7FFFFE000012099000FE3FFFB8FFE64554DF8D01E81FFEF5FCE5C3866FEC;
defparam prom_inst_10.INIT_RAM_04 = 256'h457B188F01C48FFE7CFBA024DEDFFF004000023BBFFC8799798239D23C007FFF;
defparam prom_inst_10.INIT_RAM_05 = 256'h000006EFFF41E64BF871B4CF801FFFFFFFFFFFBC100000017300003FFFFFCEF8;
defparam prom_inst_10.INIT_RAM_06 = 256'hFFFFB1000000020814000FFFFFBBFF1E953AE007C3D3FFFFFFE7C47BE1FFE800;
defparam prom_inst_10.INIT_RAM_07 = 256'h8D0793CDD8FFF9FFF1F0FFF47FFF6000000607FFF43CD908075A67009DFFFFFF;
defparam prom_inst_10.INIT_RAM_08 = 256'h0401DFFC07195B8D2F63002FFFEFFFFFFF3C80000000C205FFFFFFFFFEFFE0CC;
defparam prom_inst_10.INIT_RAM_09 = 256'hC2000000000507FFFCFFFFF7FFFC38CCAF3FD8C787FF9DFFCE6302FFFED00000;
defparam prom_inst_10.INIT_RAM_0A = 256'hC3B9BD65FF7FFF1F88487FFFF52000018E7FFFC0E3B5E0D9B9C00BFFEFFFFFEF;
defparam prom_inst_10.INIT_RAM_0B = 256'hA1DFF42E7B1899997003FF7A3F7FFF60800000000883FFFFFF613FB9FFC3C767;
defparam prom_inst_10.INIT_RAM_0C = 256'h00000002207BFFFE47B1EFFFF81F19A0BBEDFDBFFFFFDFFA140CFFFF0000008A;
defparam prom_inst_10.INIT_RAM_0D = 256'hD0D00FF9B7FFFBE075FFFFC0000043BFFFFF03C79101D860003F600FFFFFD800;
defparam prom_inst_10.INIT_RAM_0E = 256'hFFF02E38FE9878181FE07C3CFC6000000000020C3F811832223FFFFF80F8EF67;
defparam prom_inst_10.INIT_RAM_0F = 256'h00008307D08512476FFBFFFC02F77C95F9F1EDEBDC7EF8267FFBEC8003001C7F;
defparam prom_inst_10.INIT_RAM_10 = 256'hF4BFFEF1FFFF285FEFF80400404F1FF7FF04E3A07C3C3FC3E0C2033008010000;
defparam prom_inst_10.INIT_RAM_11 = 256'hF01E07E43D7038F810081F000000000000000000002C55C7FFFBFFC00F428FED;
defparam prom_inst_10.INIT_RAM_12 = 256'h000A010827141BFFFFFFFE40724184E90FFBFFFFA72BFFFFFE000056077FFFFF;
defparam prom_inst_10.INIT_RAM_13 = 256'hFEEFFFE9E607FFFFC1002CA9C7EFFFFF01F8043F21263D1000FC900000000000;
defparam prom_inst_10.INIT_RAM_14 = 256'h0FFF3CE53C4F42083F2300000000000000000F802E70FFFFFFFFFE0ED11DDFFD;
defparam prom_inst_10.INIT_RAM_15 = 256'h006F8E5CC5FFFFFFFFFFF05E6796FABF9EFF669EF3FFFFE020234A71FDEFFFF8;
defparam prom_inst_10.INIT_RAM_16 = 256'hFFE7663C9FFFE880007EF9FB9FFFFFA05FFC0B5C53F80053FFA3000000000000;
defparam prom_inst_10.INIT_RAM_17 = 256'h7F86D02CF8000FA8928000080000005E5012C003FFFFFFFFFFFF8C8DEEB5FFF9;
defparam prom_inst_10.INIT_RAM_18 = 256'hEC073CFFFFFFFFFFFFF09885EBFAFBFFFFFBAE1BFFF7A40135D9F9FA7FFFF800;
defparam prom_inst_10.INIT_RAM_19 = 256'hFEF6D7FFFFDC10031BF7F7AFFFFFE00B8114F37F800F480770000000003C61E5;
defparam prom_inst_10.INIT_RAM_1A = 256'hA7AF4FE102F0081700000092C5CCD4F803FFFFFFFFFFFFFFFF9277CF793FEFFF;
defparam prom_inst_10.INIT_RAM_1B = 256'h3FFFFFFFFFFFFFFFF3A3FB745BFBFFF5D9A6FFFFE111072CFF77EC2FDFFF01E6;
defparam prom_inst_10.INIT_RAM_1C = 256'hFEDFFFFE0441D365D45ADB1FFFC0714D1C93F880C203F9E00000333C0FFEC008;
defparam prom_inst_10.INIT_RAM_1D = 256'hB4FE003001C43480013D06E000000113FFFFFFFFFFFFFFFC717374BF7EFFFFFF;
defparam prom_inst_10.INIT_RAM_1E = 256'hFFF80DEDFFFFFFE663E6FC7FFFFFFCD97DFFFF611C266FEEA0FC9DDFF859FDB9;
defparam prom_inst_10.INIT_RAM_1F = 256'h7FFFE4C10183FF602BFD7FFF060F5A127F200945F3870001382EE0000000003F;
defparam prom_inst_10.INIT_RAM_20 = 256'hC80211FFE343F7F485D000000000000000A871FFFFFFF8CC7A9E1DFFFFFEB64B;
defparam prom_inst_10.INIT_RAM_21 = 256'h24002FFFFFFF1F03BFAABFFFFFDFFFFFFFF630A4016F900A2EFFFFC73CB6F69F;
defparam prom_inst_10.INIT_RAM_22 = 256'hFDAD1147D0777E13EFFFF0CC53FC47FA00E24FED7C07AA23C00000037D7E77F4;
defparam prom_inst_10.INIT_RAM_23 = 256'hEC07FF97FFCCA39000007A2EDAABFD31A347FFFFFFFAABF25E4FFFFFFB7BCFFF;
defparam prom_inst_10.INIT_RAM_24 = 256'h49FFFFFFFE5C7FD9C8FFFFFBFECFFFFB95620E0300E006F3BFFC66DE9071FE03;
defparam prom_inst_10.INIT_RAM_25 = 256'h10DC05805E03B0FFFF18F56EACFFE0D303FFCDFF9937C5000FD5B49C0375ED46;
defparam prom_inst_10.INIT_RAM_26 = 256'hEFD7FF7E1797803FC95EE3FFE0A69F127FFFFFFFC88F7C54BFFFFF7FBFFFDF9F;
defparam prom_inst_10.INIT_RAM_27 = 256'hFFFFFFFC53EB06B9FFFFF790FFFFEC0051C3CCF11883EFFF844306963FCB4F00;
defparam prom_inst_10.INIT_RAM_28 = 256'hF082C3C0A3BFFF834F984B1F7335E03778FFC1D7C3E87D7F18F0001CEB96FF7F;
defparam prom_inst_10.INIT_RAM_29 = 256'h5FE5C764A6FBB98FC0001BDC8B5586EFFFDFFF807F41CFBFFFFF3BBFFFFBC05D;
defparam prom_inst_10.INIT_RAM_2A = 256'hFFFFF845C159AFFFFDEE7FFFFE8C064A81DA320C933FF99D5EC50FFFC8B407F8;
defparam prom_inst_10.INIT_RAM_2B = 256'hC2E18204FBFC6F3FF283FEE00F02FF7F6DE7E06EF15D3C000006E6ACCE95F3F7;
defparam prom_inst_10.INIT_RAM_2C = 256'hA7F81FF114F40000074AE600F4B53DCFFFFE19CB6005FFFD7BD4FFFFDC110828;
defparam prom_inst_10.INIT_RAM_2D = 256'hFFDA3E84619FFFFEE7FFFFF80001FBBE80048337FC30CBB063FFD85B807FC7E1;
defparam prom_inst_10.INIT_RAM_2E = 256'h08604FFF8DA972B0FFFEB97C0F37BA47FFFFE71CF0000001ECA1CF1363197DFF;
defparam prom_inst_10.INIT_RAM_2F = 256'hFFEAC1E8000000EF16000360B47DFFFFFDC7B05017FFFFEFFFFFDD400060A780;
defparam prom_inst_10.INIT_RAM_30 = 256'hA0B12056FFFF5DFFFFFECC417ABC98200011FFCE0A23583FFF49BC17ABD387FF;
defparam prom_inst_10.INIT_RAM_31 = 256'h33FFF372076C7FFF99BB83B395F3FBFFC3A3F80000005CE8BFFFC461B7FFFFFF;
defparam prom_inst_10.INIT_RAM_32 = 256'h83E00000001850FFFFFF3721BFFFFFE610DA777FFFF60E7FFFF0022E2E841000;
defparam prom_inst_10.INIT_RAM_33 = 256'h1841E3FFFF92DFDFF0004BAB01E0200DB7F0F948763FFFF00FF5359709FFFFD1;
defparam prom_inst_10.INIT_RAM_34 = 256'hFC4ADED90FFFFE27FEB7CC79FFFF97F7E63900003DCA3FFFFFF9831FFFFFFEDA;
defparam prom_inst_10.INIT_RAM_35 = 256'h88000008FB0FFFFFFF1A8577FFFF9D4513F23FFFBF77FFFF7012E080671003FF;
defparam prom_inst_10.INIT_RAM_36 = 256'h74E7FFF9DFFFFFD00024600680003DFE23393383FFFFF17FE3E044FF7FADA7F9;
defparam prom_inst_10.INIT_RAM_37 = 256'h208140FFFFFBFFFFF20A7FFFB467FE400000079687FFFFFFF33DFFFFFFF9203D;
defparam prom_inst_10.INIT_RAM_38 = 256'h0003D7017FFFFFFF456FFFFFFF8419CDC8FFFFFFFFFFED955B10566208F7FC1B;
defparam prom_inst_10.INIT_RAM_39 = 256'h1FFFFFFFFFFDE454C19D18823FFF0C8AFF307FFFFFFFFFF9A63FFF954FFF8800;
defparam prom_inst_10.INIT_RAM_3A = 256'h087FFFFDF7FFFCF71FFFF78FFFE04000006191FFFFFFFFC4807FFFFFEB87F3DA;
defparam prom_inst_10.INIT_RAM_3B = 256'h1EC47FFFFFFFFE0DDFFFFFFC37A1B1D1FFFFFFF7FF234001A2E786FFFF862EE0;
defparam prom_inst_10.INIT_RAM_3C = 256'hFFFFFDFF1D85E3BDB1FA1FFFE3A273960FFFFFFFFFFE728FFFDC4FFFF6000000;
defparam prom_inst_10.INIT_RAM_3D = 256'hFFFFBFFFFE2EC7FFE97FFFFFA000003C3503DFFFFFFFC44BFFFFFF0178EBF67F;
defparam prom_inst_10.INIT_RAM_3E = 256'hC01FFFFFFFE3C7FFFFFFC03FD3FC0FFFF7FEFFF3008666EF6203FFF9D5275B0F;
defparam prom_inst_10.INIT_RAM_3F = 256'hFFBFFF96BDF8F3BF3FFFFC4E2CC081FFFFFFFFFF1727FFCADFFFFBE000800727;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b1;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'hFFFFFF8C71FFE1FFFFFFF8401001DCD0078EC7FFF8701FFFFFF007FFFDF9FFFF;
defparam prom_inst_11.INIT_RAM_01 = 256'hFB7FFFFF1047FFFFFC10B5DF7DAFFFFFFBFFD6AEEFF9FBDBFBFC725FF9607FFF;
defparam prom_inst_11.INIT_RAM_02 = 256'hFFF96FB7D7FFFFFFFE1AA2ABB03FFFFFFFFFE55C7FF6D7FFFFFF810001E8C801;
defparam prom_inst_11.INIT_RAM_03 = 256'hFFFA420FF15BFFFFFFFE10003AD200826CFFFFE3227FFFC81355FD3EA3FFFFFF;
defparam prom_inst_11.INIT_RAM_04 = 256'hBFFFF8EC2FFFF3007FF82E6CFFFFFF3F7F17EFFBFFFFFFFE1D2D3AAC37FFFFFF;
defparam prom_inst_11.INIT_RAM_05 = 256'h42FFFCFFFD9FFF8E4155960FFFFFFFFFF9DD1FF1F5FFFFFFFFE4001EBA40097B;
defparam prom_inst_11.INIT_RAM_06 = 256'h72CFF09D7FFFFFFF7B002F942005800FFBFE9BD9FFFFD0077E7DAF17FFFBFEFA;
defparam prom_inst_11.INIT_RAM_07 = 256'hFD84C15FFFC8006D1D37E9FFFFF1FFFFFFFEFFFFFFFFC348D839C7FFFFFFFFF8;
defparam prom_inst_11.INIT_RAM_08 = 256'hFFFFFFFFFFC73857AA41FFFFFFFFFC31E7FC639FFFFFFFFFF87BF030000003B8;
defparam prom_inst_11.INIT_RAM_09 = 256'hF8262FFFFFFFF7F432DDE6C000096E6DE02DEEFFF010087C43211FFFFCFFFBFE;
defparam prom_inst_11.INIT_RAM_0A = 256'h1F83FEF300C51F8BE7AABFFFFFFF6FFFFFFFFFFFC3199709301FFFFFFFFF90E1;
defparam prom_inst_11.INIT_RAM_0B = 256'hFFFFFFE3C975D39C3FFFFFFFFF4B505F15D1FFFFFFFFFC043FCA7000001063A0;
defparam prom_inst_11.INIT_RAM_0C = 256'h9C7FFFFFFFFF010FE63800001C80F604F20B7CC06933D74F807FFFCFFDEEF7FF;
defparam prom_inst_11.INIT_RAM_0D = 256'h07D700101E5FE9F4077FE3FFFACFFFFFFFFFF38740F7A72FFFFFFFFFD654380A;
defparam prom_inst_11.INIT_RAM_0E = 256'hFFF1C485909187FFFFFFFFC3820E85A27FFFFFFFFFBA26FB0480180A001E008D;
defparam prom_inst_11.INIT_RAM_0F = 256'hFFFFFFFFFF83BF1540002C0092E40510DAB010018FF5FFD13FDAFFCF7FA7FFFF;
defparam prom_inst_11.INIT_RAM_10 = 256'hA1000029ADE5F72FFCBFFFBFDFFFFFFFF99E05557CC2FFFFFFFDF5EF8122798E;
defparam prom_inst_11.INIT_RAM_11 = 256'h38C9F50A303FFFFFFFFC4040419942FFFFFFFFFBE3BFD94C00716044810A4837;
defparam prom_inst_11.INIT_RAM_12 = 256'hDFFFFFFF39F9888150040201061F832100000F3FFFFFA5FF0FFFFF6EBFFFFFF1;
defparam prom_inst_11.INIT_RAM_13 = 256'h0001227FB2441FBBFFE77FBFFFFF797394FFE89C0FFFFFFFF9BFB080DBB1FFFF;
defparam prom_inst_11.INIT_RAM_14 = 256'h70EB4323FFFFFFF910F81078FC1FFFEBFFFFFFCEBEDAA0220700801193200400;
defparam prom_inst_11.INIT_RAM_15 = 256'hFFFFFB0FC23C0C00650004587001C00000047C14FC9140CFFCFFEFFFFFC43ABC;
defparam prom_inst_11.INIT_RAM_16 = 256'h05FEBC3E90041FEFF7FFFFFF848FC3901259817FFFFFE7860C001376077FFF7F;
defparam prom_inst_11.INIT_RAM_17 = 256'h54601DFFFFDFE19B000D03004FEBFFFFFFFEF7390761934040803DE800000000;
defparam prom_inst_11.INIT_RAM_18 = 256'hFFFECB715C02D410380B4E000000000082BBBFFA000FFFFFFFFFFFC607AB251C;
defparam prom_inst_11.INIT_RAM_19 = 256'hF2621FC003FFEEF7FFFF0502C70DFFE90800FFFFFDF88FC006E0C012FBFFFFFF;
defparam prom_inst_11.INIT_RAM_1A = 256'h03FFFBFDEC7A40018B2079F7BEFFFFFFFF0BEF3103F5A186039F880000000030;
defparam prom_inst_11.INIT_RAM_1B = 256'hF89CF4B2FE0632074A400400000003DB6AAD3DD8FFFFFFFFFF8378077137A267;
defparam prom_inst_11.INIT_RAM_1C = 256'hA33F861FFBFF87FFC0E073BB02705DE0BFFFFDE038D0019C38206E5FFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1D = 256'hFEEFFE094C00E6AE08679EFFFFFFFFFE3B8FF6078188036EB00000000000DE00;
defparam prom_inst_11.INIT_RAM_1E = 256'hF53EA00F000EC04C00000000005AF2895BC007FFFBFFFFE0C03BE79D5AEB380B;
defparam prom_inst_11.INIT_RAM_1F = 256'hA803FFFFFFFFF0E00FF85C824A4F06069F8C06560034368279FE9FFE7DF7FFEF;
defparam prom_inst_11.INIT_RAM_20 = 256'h600315001D37A0001DCBF99F7FF7FFFCBAE280004DFF4F00000000000F2BD270;
defparam prom_inst_11.INIT_RAM_21 = 256'h99D1B369F327800000000802ED51D40D00FFFFFFFFF078228A66258259E019C6;
defparam prom_inst_11.INIT_RAM_22 = 256'h3FFFFFDFFC3011A60093670A70500E6200E6C00CA6F00027E0A093F17FFFFF19;
defparam prom_inst_11.INIT_RAM_23 = 256'h2DA00778BC0001700000030FFFFF819CA992B8FE1AC000000004187F6DDF585C;
defparam prom_inst_11.INIT_RAM_24 = 256'hABCE34017000000000C61F855781A200FFFFEFFF1D045CCECD8C5C9C00040000;
defparam prom_inst_11.INIT_RAM_25 = 256'hFFFFFF4768723EBB783053000860041ED8019AAC00020440000000002000722B;
defparam prom_inst_11.INIT_RAM_26 = 256'h00E497C0400E8000000000000B46856392404EB4000000014987F4B04706603F;
defparam prom_inst_11.INIT_RAM_27 = 256'h8321FE000004000413D5581940B6DFFFFFFFE3DA771FBB083075C00000000464;
defparam prom_inst_11.INIT_RAM_28 = 256'hFED1DA39BFAA5862916800008201DB00780DE00000008000000908DB45D92D1D;
defparam prom_inst_11.INIT_RAM_29 = 256'hB2780001000000002FBFD48FC4C1A3678BFF80004080110D3DBE6B2AA2D8FFFF;
defparam prom_inst_11.INIT_RAM_2A = 256'h7F2000001159E3FFF91E852033FFFFFFF8F3ECAFEA0802A04E000020008E807C;
defparam prom_inst_11.INIT_RAM_2B = 256'h7B0DEFF573059297800000002B600F5F9C0000002000001FFC52C01B78C54D74;
defparam prom_inst_11.INIT_RAM_2C = 256'h801000000001FF41EA60092AF1F939FFE8004008678FFFECCF02F0347FFFFFF8;
defparam prom_inst_11.INIT_RAM_2D = 256'h0002013C6BFBDFD541AC5C3FFBFFFF8CD5AB7F0F47E144E000000008D40F9A47;
defparam prom_inst_11.INIT_RAM_2E = 256'hCFFE5C032F657C00000003DC03EC99E80080000000FF45D34C01024DFF03FFFF;
defparam prom_inst_11.INIT_RAM_2F = 256'h20000025FF43D847E000FB1801FFFFE101CFFF7E5EFFFE84500D87FFFFFF06F2;
defparam prom_inst_11.INIT_RAM_30 = 256'h33FFFEFFDFFFD9800FE97FFFFFE3D120D1CEE0C1428F00000001331BF2D47E40;
defparam prom_inst_11.INIT_RAM_31 = 256'h79B0E4A42720000000DC897CE71F80000000097FC39E6DF6C053A4002FFFFC90;
defparam prom_inst_11.INIT_RAM_32 = 256'h003C7F039A1ACFEA3F1D0007FFFFC83F7FFFFFFFFFEF2005E29FFFFFC32A2185;
defparam prom_inst_11.INIT_RAM_33 = 256'hFFFFFFFFFFF400723FFFFFC0A164625DD8F1BE79F00000001DE2FE20CFE10040;
defparam prom_inst_11.INIT_RAM_34 = 256'h75C9C47E00000023FB3F95A3FC01000001FFC38F809FA208A1F8003FFFE9D63F;
defparam prom_inst_11.INIT_RAM_35 = 256'hFFC1CDA50ED960B9F8000FFFFF9FDFBFFFF7FFFF0F801581FFFFA56F89CFD9CC;
defparam prom_inst_11.INIT_RAM_36 = 256'hFFFFF7F91C3FC47FFFE1A7BC87889DFF90563F0000000277FFE0A9FF00000009;
defparam prom_inst_11.INIT_RAM_37 = 256'hFF8FC0000003B9FFF9EC6FF00000007FF0E69D9B4CD8124F8002FFFFC77FFFEF;
defparam prom_inst_11.INIT_RAM_38 = 256'h615AE414B10AEDF00127FFF3FFF3FFFFFFFFDF6EFBC46FBFC03312C921903D11;
defparam prom_inst_11.INIT_RAM_39 = 256'hFFBFF704EB09ABC0B6A9A008231EBC9F67F000000045FFF853CFF400006147F4;
defparam prom_inst_11.INIT_RAM_3A = 256'hF84000003D5F7E1043EE0000082FF819A3CD3FD4432E8E0007FFFE7BFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3B = 256'h2706EA9875CFF000EFFFFFFFFFFFFFFFFFFF7040C047A0D23E3620008BB8EF33;
defparam prom_inst_11.INIT_RAM_3C = 256'hFFF0E4D019001485AB20B503F6EE08FE0000007D1FFF8D58FBC4001045FE1CD7;
defparam prom_inst_11.INIT_RAM_3D = 256'h00085EDFFF218E3EF0480471FB0E4953405539EA23EE001BFFFEFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3E = 256'h3E18CE8A6880037FFFFFFFFFFFFFFFFFFFC5EE05803DF1F6A166207CCB4E1F80;
defparam prom_inst_11.INIT_RAM_3F = 256'hFFFF000015FFBD7E0C403D71831FFC000001A4FFF8E50FFDC0127FFE87759438;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b1;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'h0000000931EDFFFFFFFFFFFFFFFFBFFFFFFF679FFFFFFFFFFFFFFFFFFFFFF404;
defparam prom_inst_12.INIT_RAM_01 = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFB004401ABBFFFFF3FFFFFFFFFFFFFFB800000;
defparam prom_inst_12.INIT_RAM_02 = 256'h683F37FCD7FDFFFFFFFFFFF600000000000000403F7EFFFF767FFDFF87DBFFFF;
defparam prom_inst_12.INIT_RAM_03 = 256'h000021597FFFFFFFFFFFFCFFBA7FFFFFDC6DBFFFFFFFFFFFFFFFFFFFFFC00012;
defparam prom_inst_12.INIT_RAM_04 = 256'hE7DDD7FFFFFFFFFFFFFFFFFFFE84081B3F91FDFFFFFFFFFFFFFFFE1000005000;
defparam prom_inst_12.INIT_RAM_05 = 256'h7FFECFFFFFFFFFFFFFFEC000005F0000000001397DFFF9FFFFFFC819F61D8007;
defparam prom_inst_12.INIT_RAM_06 = 256'h0000184EF7FE79FFFF300210006001999A76FFFFFFFFFFFFFFFFFFFF880045FE;
defparam prom_inst_12.INIT_RAM_07 = 256'hE0FCFFFFFFFFFFFFFFFFFFFC00037FFFFFBBFFFFFFFFFFFFFED000003FF00000;
defparam prom_inst_12.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFBE4000002FFF60000000021B79DFFFFF4C0208100108032B43;
defparam prom_inst_12.INIT_RAM_09 = 256'h0100637FB41E8600000040400B664A2D02CFFFFFFFFFFFFFFFFFFF8024FDFFFD;
defparam prom_inst_12.INIT_RAM_0A = 256'hBFFFFFFFFFFFFFFFFFFFE008FFFFEFFFFFFFFFFFFFFFB20800004FFFFC000000;
defparam prom_inst_12.INIT_RAM_0B = 256'hFFFFFFFFFFEF42000017FFFF400000005818FFE807A0800008205002C86A8860;
defparam prom_inst_12.INIT_RAM_0C = 256'h01FF8696003008200000001049C0027FFFFFFFFFFFFFFFFFFFFC073EFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFF203BFFFFFFFFFFFFFFFFFFFF74000001FFFFD300000000;
defparam prom_inst_12.INIT_RAM_0E = 256'hFFFFFFFFFB000005DFFFABE0000108007FE020800C0100000000001A800037FF;
defparam prom_inst_12.INIT_RAM_0F = 256'hFE068000000200000000184E081FFFFFFFFFFFFFFFFFFFFFF0AFBBBFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFE83FDFFFFFFFFFFFFFFFFFFEF340000F7FFF05F2000000241F;
defparam prom_inst_12.INIT_RAM_11 = 256'hFFFFFD008003EFAF93FF7000100539F786440C000000002000038AEF0DFCFFFF;
defparam prom_inst_12.INIT_RAM_12 = 256'h910300000000000000622DC1FFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_13 = 256'hFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFBB40400FFFFFA47FF6A04100CFFBE1;
defparam prom_inst_12.INIT_RAM_14 = 256'hFFA4000FFFE5997FFFE007F9FE7FDB837000000000001080009D1C73FFFFFFFF;
defparam prom_inst_12.INIT_RAM_15 = 256'h10000C000008000001844F5FFFFFFFFFFFFFFFFFFFF43EFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_16 = 256'hFFFFFFFFFDFB7FFFFFFFFFFFFFFFFFFFFE000DFFFED6FFFFE93FF7DFFFFDF962;
defparam prom_inst_12.INIT_RAM_17 = 256'h8002FFFFF57FFFE51FFFFFFFFEEFF88000F000000000000042EC5FEFFFEFEFFF;
defparam prom_inst_12.INIT_RAM_18 = 256'h0240018100000000F8FFFDFFFFEFFFFFFFFFFFFF7FFFBFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_12.INIT_RAM_19 = 256'hFFFFFFFFFFFFEFFFFFFFFFFFFFFFFB68047FFFDDBFFFFE3DFFFFFFEFFF7A0000;
defparam prom_inst_12.INIT_RAM_1A = 256'hFFFFF5B7FFF2FFDFFFEFFFFFE6C00000000068400000602233FFFFBFFFBFFFFF;
defparam prom_inst_12.INIT_RAM_1B = 256'h0000800000003D3FDAFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFEC400;
defparam prom_inst_12.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFBF127E77FEEBF79FA3FFCFDFFFFFFFE60000000;
defparam prom_inst_12.INIT_RAM_1D = 256'hF29FEFA97FFFCBFFFFFFFFE00000000101010000000B0EFFCFFFFFFF7FFFFFFF;
defparam prom_inst_12.INIT_RAM_1E = 256'hC0A0000002C3FFDFDFEFFFDFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFEB60BCF7;
defparam prom_inst_12.INIT_RAM_1F = 256'hFFBFFFFFFFFFFFFFFFFFFFFBF1BFA7735FFF3FBFFFFCFFFFFFFFF8000000FF01;
defparam prom_inst_12.INIT_RAM_20 = 256'hFFFBFFFFFEBFFFFFFF7618000BFE51400055002020FFAFFFF7FFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_21 = 256'h0100004F97DFFFFFFFFF7FFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFEFFCBFFB7F4F;
defparam prom_inst_12.INIT_RAM_22 = 256'hFBFFFFFFFFFFFFFFFFFFBFFFFFBE9FFFFCDEFFFFC7FFFFFFF4800005E2238200;
defparam prom_inst_12.INIT_RAM_23 = 256'hD4EFFFD5FFFFFFF6400001C084BC000025010307FBFFFBFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_24 = 256'h40016FDFDBFFFFFFFBFFFFFFFFFF7F7FFFFFFFFFFFFFFFFFFFFBFFFFFBA7FFFC;
defparam prom_inst_12.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFF3CFFFFF967FFECF2EFFABFFFFFFFF400003E31A21800000;
defparam prom_inst_12.INIT_RAM_26 = 256'hEFF7FFFFFFFE480003E028FDE00000100269F7F9FBFDFFEFFFF7FFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_27 = 256'h000FFDFFF77B3FE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCC7FFFD1967FEEDF2;
defparam prom_inst_12.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFECFFFF96077E34FFAC36F7FFFFFFF0002074B2C98E00000400;
defparam prom_inst_12.INIT_RAM_29 = 256'hFDFFFFFFFC8000363AFDCAE0000000000EDFFFBCFCD97FFFFFFFFFFFDFFFFFFF;
defparam prom_inst_12.INIT_RAM_2A = 256'h87FFFF3F33DFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFECFFE9DFCE1DAFFF778;
defparam prom_inst_12.INIT_RAM_2B = 256'hFFFFFFFFFFFF557E09FFCA0AFFFF34FF7FFFFFFD20001CC7E80FFE0000000003;
defparam prom_inst_12.INIT_RAM_2C = 256'hFFFFFFA00007D827733F90000000001EEFFE7FF7B9FFFBFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2D = 256'hF3FFFFBFEEDFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFDB45FFFFF97FFFECBFFF;
defparam prom_inst_12.INIT_RAM_2E = 256'hFFFFFFFFFFFD06FFFF394FFFF40FFBFFFFFFD60043EB3EC637FC00000000003C;
defparam prom_inst_12.INIT_RAM_2F = 256'hFFE60200FD4E40881F00000000000C3E7FDBDDFBF1FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_30 = 256'hB7FEFFEEFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFED8FFFF8CE3FFF8BFFC7FFF;
defparam prom_inst_12.INIT_RAM_31 = 256'hFFFFFFEFE37FFFC8DB3FFA16FF5FFFFFFD40003F29401051F00000000000BF3F;
defparam prom_inst_12.INIT_RAM_32 = 256'hD0203FE4400165FD00005880001FCFFFE6BEFBDFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_33 = 256'h9EFE7FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE2FFFF299BBFEEFFF61FFFFFF;
defparam prom_inst_12.INIT_RAM_34 = 256'hFFFE7FAF7FD44E5B3D8FFFB005FFFFF800017C5802B9C780001DEA01004DFFFB;
defparam prom_inst_12.INIT_RAM_35 = 256'h0017AF351FB5F80008001080C3EEF597FCFFFEFFFBFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_36 = 256'h6167FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEB7F30FF1B6136FF2007FFFFFC0;
defparam prom_inst_12.INIT_RAM_37 = 256'hFFFCEF78A7FE135DDAD14007FFFFF00047E6E501E79E000580062433F8BFE3FE;
defparam prom_inst_12.INIT_RAM_38 = 256'hFCCE325FFBA00026020026DCFDFBF7FCDF7FFBFFFF7FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_39 = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFE7E7C708FFFFC20FEF9F000FFFDDC284F;
defparam prom_inst_12.INIT_RAM_3A = 256'hDFD793DFFE1BDFFCF4001FFFFF5D73FFA0EFDCBF780000002001A37FFF4FFFAF;
defparam prom_inst_12.INIT_RAM_3B = 256'hE5FF5F5F000000002037FFEFE77FA7E76B3FFFFFFFFFFFFFFFFFFFFFFFFFFFA7;
defparam prom_inst_12.INIT_RAM_3C = 256'hFDFFFFFFFFFFFFFFFFFFFFFFFFFFFD73FD2BFFBF827FFD7E8007FFFFFFDDFFF5;
defparam prom_inst_12.INIT_RAM_3D = 256'hC88FFFF4DFFFFF3B00FFFFFFFFFFFE5CBF387FF00000000058CCFFFE19E76E1B;
defparam prom_inst_12.INIT_RAM_3E = 256'hD6FEFC0000000026333FFF9E79D9E3FF7FFFFFFFFFFFFFFFFFFFFFFFFFFE967F;
defparam prom_inst_12.INIT_RAM_3F = 256'hFF7FFFFFFFFFFFFFFFFFFFFFFFF427FCAFFFC04BBC1FFF007FFFFFFFFFFFCD77;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b1;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'h3FE3F0FF2FF3F03FFFFFFFCEFFFCB2FFF4E7C00000800B40FEF5F87E4423314F;
defparam prom_inst_13.INIT_RAM_01 = 256'hFCF00000000037FEFFBFE7E3F93D77FFFFFFFFFFFFFFFFFFFFFFFFFFCB8AFE98;
defparam prom_inst_13.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFBE5EFBD8BC8947E17FEFE07FFFFF9A765FF8A5CF9;
defparam prom_inst_13.INIT_RAM_03 = 256'h1F5ECCFE3F83FFFFFCEFCDAFF1B9FB9FAF0000000004FF9FEB79F167BEFF6FFF;
defparam prom_inst_13.INIT_RAM_04 = 256'hE0000000848EBDFFFFF03877DFDFFFFFFFFFFFFFFFFFFFFFFFFFFEFEAFFFFAB0;
defparam prom_inst_13.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFDFD6FD67ACBFD70E7F27E0BFFFF289C58F7F2633E2F9;
defparam prom_inst_13.INIT_RAM_06 = 256'hE39F08F83FFFF09632D0EF8487DDF6BE00000002236F779F7B873FF9FFFFBFFF;
defparam prom_inst_13.INIT_RAM_07 = 256'h000000015FFFDEFE40817EFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFDFDE4FB23F2;
defparam prom_inst_13.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFDFFBBFA4BCFFFB1F7B53C0FFFF9D117E4DDCC84FBDD87E0;
defparam prom_inst_13.INIT_RAM_09 = 256'hDC4E07FFF9DB6C45D7671097FFFEFC000000003FFDFFFFF967FFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0A = 256'h000C3FFFFFFFE6187FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FE61C780FFF1DF9;
defparam prom_inst_13.INIT_RAM_0B = 256'hFFFFFFFC7FFFFE0BF3F2920FFFEFFE5213807FF0BDFBE06CE2B2B3F777BF8000;
defparam prom_inst_13.INIT_RAM_0C = 256'hC05FF85486C0E96AD4564757E7F02000002DFFFFF8E011F978DEF7FFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0D = 256'h13FFDF9E7F1AED1FFF7DFFFFFFFFFFFFFFCFFFFFFFFF831BFF2C01BFE37F9264;
defparam prom_inst_13.INIT_RAM_0E = 256'hBEFE7BFFFFE0C3BFEB81EFF91FE6B16017FC280D73F288B54BCB2C5F7F400100;
defparam prom_inst_13.INIT_RAM_0F = 256'hFE1DFC6001D3AE3971371FEFF00000009FF7FFDF9F78A7EFFFDFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_10 = 256'hDFFFFDE7A0F8DDFFFFFFFFFFFFFFFFEF7FD03F3BF83E3BFC787BF207E55CD803;
defparam prom_inst_13.INIT_RAM_11 = 256'hE81FFC7E0BE6FFBB087FEBF85F20017F0CA9207E0CCCB82C3E7F6CFFFB0003DF;
defparam prom_inst_13.INIT_RAM_12 = 256'hD8107FF842BE8584BCAF9FFE4200FFF4FFFEFFF90F375FFFFFFFFFFFFFFFF38F;
defparam prom_inst_13.INIT_RAM_13 = 256'hFFFFF3847F7DFFFFFFFFFFFFFFFD01FEE7EC1F83E5DFE2BF1DBCFD8F86005FC2;
defparam prom_inst_13.INIT_RAM_14 = 256'hFCC7E05ECBFBEFD5DE3CB1D1E00FE1E1687FFF8DB6E0B0DCF6143FD023CFDEFE;
defparam prom_inst_13.INIT_RAM_15 = 256'h3FFFF8AED20E1EBCFFA34ECCF3F7FFFFFFE69118FEFFFFFFFFFFFFFF37C07F50;
defparam prom_inst_13.INIT_RAM_16 = 256'hF932481FFFF7FFFFFFFFFF9E5D1FF8FF71E0170D7EF84C4FB75EB23803F85938;
defparam prom_inst_13.INIT_RAM_17 = 256'h7A01E12B8EC74FE65F22E700F832FB3FFFFF94238103F8605004333EFFFEDFF3;
defparam prom_inst_13.INIT_RAM_18 = 256'hFFF291B0663E509FFFDDFFFF35F9FCFEEFBCEFFFFFFFFFFFFFFFEFBF45FF2F91;
defparam prom_inst_13.INIT_RAM_19 = 256'h707BFFFE7FFFFFFFFFFE85E13FC3C1BC007078F5E9BFFC37FA3BC0180E324FFF;
defparam prom_inst_13.INIT_RAM_1A = 256'h6A0789ED9BFFCFF2B8F8040286E1FFFFFE5F8C86CEE01E301E1FFCFBFBFFF859;
defparam prom_inst_13.INIT_RAM_1B = 256'hC904B898F01EB00173FFFEF7FFDE7E603FEFFF4BFFFFFFFFFE803C0A80D13E00;
defparam prom_inst_13.INIT_RAM_1C = 256'hFBDFCFFFFFFFFFFF8070038CA91F01F106FE3FD8FFD3FD8E3E00009618FFFFFF;
defparam prom_inst_13.INIT_RAM_1D = 256'h87E5FEFFCAFE070F000025263FFFFFF1CA6F1B1C1F94FE0E3FBEDFF7E1FBBA82;
defparam prom_inst_13.INIT_RAM_1E = 256'hB9E760F7FDFFF2DFFFBBFC99DE975030F7FFFFFFFFFFFFE90798706F0BC078FC;
defparam prom_inst_13.INIT_RAM_1F = 256'hFD1FFFFFFFFFFFFE78017E3BC07C7739F27B6FE17F020780000EE40FFFFFFE57;
defparam prom_inst_13.INIT_RAM_20 = 256'h6FEFF3CFF003E001034401FFFFFF936C7CA55F91FFFB1FFFFFEFFBFF9F4F1877;
defparam prom_inst_13.INIT_RAM_21 = 256'h164BC1FFFFA3DFFFBEDFF887D98BFFFF7EFFFFFFFFFFFE84000FFEA01F0E263F;
defparam prom_inst_13.INIT_RAM_22 = 256'hFFFFFFFFFFFFCC001FFFA40F83C71FF67EF36BEF00F00000438CFFFFFFC4369F;
defparam prom_inst_13.INIT_RAM_23 = 256'h1C7CCFE03C0004170F1FFFFFF30B67E2EAB1FFFFFC33FFFDBFFE21E608FFFFC6;
defparam prom_inst_13.INIT_RAM_24 = 256'h5CFFF7FF96FFFFE7FF85FDE8F03FF1FFFFFFFFFFFFF8001FFFEC07E0FFE9FF2F;
defparam prom_inst_13.INIT_RAM_25 = 256'hFEFFFFFFBFB007FF7783F03FFDFC32D27E29F01F8004029D23FFFFFCA3D9F8A4;
defparam prom_inst_13.INIT_RAM_26 = 256'hABFC1FC00660A5B4FFFFFE590E7F2A203FFFF7C1CFFFFFFFFFFE0E134DFC1BFF;
defparam prom_inst_13.INIT_RAM_27 = 256'hFFFDFE33FFFDFFF79FE7A1FDFF8FFFFFFFFFFFF7D81BF03E85F80BFFFF2FB4BF;
defparam prom_inst_13.INIT_RAM_28 = 256'hFFFFFFFF99C78709FC00FFFDFFFD7FE0FE07E001F830BF1FFFFF182EBFC8C94F;
defparam prom_inst_13.INIT_RAM_29 = 256'h83F8000F051AE7FFFF8BE4CFE2A62BFFFF7F877FFFFFF5E998082FFFD3DFFFFF;
defparam prom_inst_13.INIT_RAM_2A = 256'hF3E1DFFFFFA11C6633075FF13FFFFFFFFFFBFFFE1FDC00FF000FC790FF0FFA3F;
defparam prom_inst_13.INIT_RAM_2B = 256'hBFDFFC5EE6800E0003C06B7FFFFC1F01FC000DC0902C7FFFCDE563F8AC88FFFF;
defparam prom_inst_13.INIT_RAM_2C = 256'h0003F832269FFF85354BFF29E39FFFFDF84FFFFFFE68FF4468D1FC5FDFFFFFFF;
defparam prom_inst_13.INIT_RAM_2D = 256'h3CFFFFFFF8F6B541EE7F07EFFFFFFFFEBBCF0EBA0008000000006FFE7F4680FF;
defparam prom_inst_13.INIT_RAM_2E = 256'h0406C076C0040000000CDEFF7980FF8003FF85D563FF8BB704FFCC0963FFFFEE;
defparam prom_inst_13.INIT_RAM_2F = 256'hFFE09CF41E043E127FF1017CFFFF7B851FFFFFBE3B6B7879FFC4DFFFFFFFFFFC;
defparam prom_inst_13.INIT_RAM_30 = 256'hFFF9FFFA758281F7F0F7FBFFFEFFBA800373107C3FF00000021FFF8F807FC000;
defparam prom_inst_13.INIT_RAM_31 = 256'hDE1D0E0FFF0000401A7D9F803FF0002FFC3C1080313D613FFC59CF1FFFFEC32F;
defparam prom_inst_13.INIT_RAM_32 = 256'h8529819C0A709FFF9933F1FFFD8169FFFFFF7D7E07D637FC2FFFFFEFFFFA0001;
defparam prom_inst_13.INIT_RAM_33 = 256'hFFBE1F2DFE45FF01DFFFBEFFFFA800573C078C0FC00FFC03ADE7E03FC0001FFF;
defparam prom_inst_13.INIT_RAM_34 = 256'h3F0280F01FFFF83849C07FF0001FFFF1947660CE174FFFE2DCEF3FFF806A7FFF;
defparam prom_inst_13.INIT_RAM_35 = 256'h76896C274FFFF8A78CE5FD80148FFFFFF87F119D97FFC17FFFFFFFFE8C0001C7;
defparam prom_inst_13.INIT_RAM_36 = 256'hFE438EE9BFF027FFFFF6AED00001FB3401801C07FFFF00B6007FF80019FFFC3E;
defparam prom_inst_13.INIT_RAM_37 = 256'h7B8F07FFFFF018E1FFFC00067FFF4748765A50CFFFFF34B19EFF003A03FFFF9F;
defparam prom_inst_13.INIT_RAM_38 = 256'h2582C7FFFFC4B603F0003C48FFFFFF1FBD690BFFFE34FFFBF7EBA800028FF080;
defparam prom_inst_13.INIT_RAM_39 = 256'h0C423F3F077FFFFFFFF40000795820347183FFFFFFFC8FFFFC00077FFFF8AF60;
defparam prom_inst_13.INIT_RAM_3A = 256'h70FFFFFFFC01FFF00001FFFFFF193492428FFFFFF99E201FEB7FC63FFFFFFFE7;
defparam prom_inst_13.INIT_RAM_3B = 256'h9FFFFBFE35C9C47FFC608FFFFFFFFFC110CFFFC2FFFFFFFFE90000181B00044C;
defparam prom_inst_13.INIT_RAM_3C = 256'h0AFFF0BEEFFFFDDA00000721C00291387FFF182000162000007FFFFFF0DF8D55;
defparam prom_inst_13.INIT_RAM_3D = 256'hF5040000000000003BFFFFFF0D8DFF1FFFFFFFC6AADA0C4300A3FFFFFFE18E50;
defparam prom_inst_13.INIT_RAM_3E = 256'hFF8BF895FA3F1180ECFFFFBBF0BE4100D7FC5FFFFFFFFE200003DC3005D6CE1F;
defparam prom_inst_13.INIT_RAM_3F = 256'hFF395FFFFEF9A80001F10787D5B39FE8000000000000001FFFFFFFF87F01DFFF;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b1;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'h0000000000001FFFFFFFFF000F87FFFFBAFF3902AFF046DF3FFFEFFDBE28401F;
defparam prom_inst_14.INIT_RAM_01 = 256'hFFC72F7A0DA67F8FFFFFBE7C67EC2FFFC27FFFBFFFF000007C2CF0070887F800;
defparam prom_inst_14.INIT_RAM_02 = 256'hF8FFFEFF1000003F852F005661FC000000000000004FFFFFFFFFFF0003FFFDE7;
defparam prom_inst_14.INIT_RAM_03 = 256'h0000000001FFFFFFFFFFFF01FFFFB8FFF8773F3F88FFE7FFFEF5FCE5C3866FF3;
defparam prom_inst_14.INIT_RAM_04 = 256'h8655A98EFFFD7FFE7CFBA024DEDFFCFFBFFFFDC4400007E185E773B1FC000000;
defparam prom_inst_14.INIT_RAM_05 = 256'hFFFFF9100001F87208888C3F8000000000000043EFFFFFFFFFFFFFFFFFFFCEFF;
defparam prom_inst_14.INIT_RAM_06 = 256'h00004EFFFFFFFFFFFFFFFFFFFFBBFFE0E64D177FEB8FFFFFFFE7C47BE1FF17FF;
defparam prom_inst_14.INIT_RAM_07 = 256'h11AEFFFFD7FFF9FFF1F0FFF47FC09FFFFFF9F800003F1E1DD3C61F0000000000;
defparam prom_inst_14.INIT_RAM_08 = 256'hFBFE200007E19234631F00000010000000C37FFFFFFFFFFFFFFFFFFFFEFFFF0F;
defparam prom_inst_14.INIT_RAM_09 = 256'h3DFFFFFFFFFFFFFFFFFFFFF7FFFFC0F0C95FABFEFFFF9DFFCE6302FFF12FFFFF;
defparam prom_inst_14.INIT_RAM_0A = 256'h83C3B74FFF7FFF1F88487FFC0ADFFFFE71800000FC3A054787C0000010000010;
defparam prom_inst_14.INIT_RAM_0B = 256'h5E20002F83BB8787F0000085C080009F7FFFFFFFFFFFFFFFFFFFFFB9FFFC0786;
defparam prom_inst_14.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFF8E7EFFFFFE01E2E3BE3E8FFFFFFDFFA140CFF00FFFFFF75;
defparam prom_inst_14.INIT_RAM_0D = 256'hD9DEBFF9B7FFFBE075FFC03FFFFFBC40000003F81EFFC7E000009FF0000027FF;
defparam prom_inst_14.INIT_RAM_0E = 256'h00002FC0FE87F818001F83C3039FFFFFFFFFFFFFFFFFFFC1CEFFFFFFFF00F5D7;
defparam prom_inst_14.INIT_RAM_0F = 256'hFFFFFFFFFFFFE19F5FFBFFFFFD063ABBF9E7EDEBDC7EF8267FF0137FFCFFE380;
defparam prom_inst_14.INIT_RAM_10 = 256'hFEFFFEF1FFFF285FFC07FBFFBFB0E0000004FC0003FC3FC01F3DFCCFF7FEFFFF;
defparam prom_inst_14.INIT_RAM_11 = 256'h001FF81BFEFFF807EFF7E0FFFFFFFFFFFFFFFFFFFFCEFF7FFFFBFFFFF06A4FFB;
defparam prom_inst_14.INIT_RAM_12 = 256'hFFFFFFFFB64487FFFFFFFFFF8559B4FF5FFBFFFFA72BFFFF01FFFFA9F8800000;
defparam prom_inst_14.INIT_RAM_13 = 256'hFEEFFFE9E607FFC03EFFD3563810000001FFFBFF1C5E02EFFF036FFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_14 = 256'h0FFFFFF6E3C0BDF7C0DCFFFFFFFFFFFFFFFFF16C5E0FFFFFFFFFFFF0A33BCFFB;
defparam prom_inst_14.INIT_RAM_15 = 256'hFF87E0C33FFFFFFFFFFFFF94679CFA7F9EFF669EF3FFF01FDFDCB58E02100000;
defparam prom_inst_14.INIT_RAM_16 = 256'hFFE7663C9FFC177FFF810604600000005FFFD4D83007FFAC005CFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_17 = 256'h7FEF39E407FFF0030D7FFFF7FFFFFFA2B7E63FFFFFFFFFFFFFFFF1C5F277EFF9;
defparam prom_inst_14.INIT_RAM_18 = 256'hA3FFFFFFFFFFFFFFFFFF318EEFF9FBFFFFFBAE1BFF085BFECA26060580000000;
defparam prom_inst_14.INIT_RAM_19 = 256'hFEF6D7FFC023EFFCE40808500000000BF980F9007FF037FD0FFFFFFFFFC01DA6;
defparam prom_inst_14.INIT_RAM_1A = 256'hADD1C01EFD7FF7E8FFFFFF6D0FA04C07FFFFFFFFFFFFFFFFFFE717CE7D7FEFFF;
defparam prom_inst_14.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFC8FFF7BC7FBFFF5D9A6FFF01EEEF8D300881010200001F9;
defparam prom_inst_14.INIT_RAM_1C = 256'hFEDFFC01FBBE2C9A2BA520E000007C912C30077F0DFC071FFFFFCC4FA0013FFF;
defparam prom_inst_14.INIT_RAM_1D = 256'h6C01FFC7FE3BF37FFEC0B19FFFFFFFFFFFFFFFFFFFFFFFFF94FBFBBCFEFFFFFF;
defparam prom_inst_14.INIT_RAM_1E = 256'hFFFFF21FFFFFFFFAD3E5BC9FFFFFFCD97DFF001EE3D990115F026220005EB61A;
defparam prom_inst_14.INIT_RAM_1F = 256'h7FC01B3EFE7C009FD40280000787290600DFF2BA0C7EFFFEC2F61FFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_20 = 256'h37FC6E001DBC0803342FFFFFFFFFFFFFFF4A46FFFFFFFF5A78BFF3FFFFFEB64B;
defparam prom_inst_14.INIT_RAM_21 = 256'hA3FFFFFFFFFFEBCDF81F7FFFFFDFFFFFF009CF5BFE906FF5D1000007DAA3B580;
defparam prom_inst_14.INIT_RAM_22 = 256'h0252EEB82F8881EC100000F65ECEC005FF5DB012E3F845683FFFFFFC9D8B5006;
defparam prom_inst_14.INIT_RAM_23 = 256'h0FF800700013F06FFFFF83606CCC0088D06FFFFFFFFC7BF3FF7FFFFFFB7BCFFC;
defparam prom_inst_14.INIT_RAM_24 = 256'h17FFFFFFFF8F7C7EAFFFFFFBFECFFF046A9DF1FCFF1FF90C40007A5C2F3001FC;
defparam prom_inst_14.INIT_RAM_25 = 256'hEF23FA7FA1FC4F00001E9D011C001F2BFC00380007D03AFFF0561D4C0381F495;
defparam prom_inst_14.INIT_RAM_26 = 256'h102E003430687FC0B095E00002CF3D10FFFFFFFFF2EFFD8F7FFFFF7FBFFFC060;
defparam prom_inst_14.INIT_RAM_27 = 256'hFFFFFFFF1FFBDF27FFFFF790FFF013FFAE3C330EE77C100007B6D9CE0034B0FF;
defparam prom_inst_14.INIT_RAM_28 = 256'h0F7D3C3F5C4000039E4667008CCA2FC8868028303C17818FB80FFFE14F313D6F;
defparam prom_inst_14.INIT_RAM_29 = 256'h403BA09B590356803FFFE5F9D771B6AFFFDFFFEBFEB77CFFFFFF3BBFFC043FA2;
defparam prom_inst_14.INIT_RAM_2A = 256'hFFFFFD77BF979FFFFDEE7FFF0173F9B57E25CDF36CC001ED541300003747F807;
defparam prom_inst_14.INIT_RAM_2B = 256'h3D1E7DFB0400710A0980011FF07D00802FA01F9102AF03FFFFFB8E99D6F107F7;
defparam prom_inst_14.INIT_RAM_2C = 256'hE007E000C80BFFFFF943FA1BEC896DCFFFFFAFFFAFD3FFFD7BD4FFC023EEF7D7;
defparam prom_inst_14.INIT_RAM_2D = 256'hFFE5FF37BF7FFFFEE7FFF007FFFE04417FFB7CC8003CF4C5E00027A43F80503F;
defparam prom_inst_14.INIT_RAM_2E = 256'hF79FB0000ED3C27000014683F0F033A0000000240FFFFFFE2CE80FB080037DFF;
defparam prom_inst_14.INIT_RAM_2F = 256'h0009A817FFFFFF2131FFFC7032FDFFFFFEBE7F7BEFFFFFEFFFFC22BFFF9F587F;
defparam prom_inst_14.INIT_RAM_30 = 256'hDFFFD7B9FFFF5DFFFF0133BE854367DFFFEE000F16C3380000B6406860152000;
defparam prom_inst_14.INIT_RAM_31 = 256'hCC0003AB7FDC000066443C60135004000CD007FFFFFF8B07FFFFF95917FFFFFF;
defparam prom_inst_14.INIT_RAM_32 = 256'hD01FFFFFFFE807FFFFFFC1213FFFFFFBFF09903FFFF60E7FC00FFDD1D17BEFFF;
defparam prom_inst_14.INIT_RAM_33 = 256'h679807FFFF92DFF00FFFB454FE1FDFF24800CED3AE00000FF005EC185800001E;
defparam prom_inst_14.INIT_RAM_34 = 256'h007CC217000001D8001C0E280000181019C6FFFFC001FFFFFFFE989FFFFFFF77;
defparam prom_inst_14.INIT_RAM_35 = 256'h77FFFFF262FFFFFFFFEE85F7FFFFEEFAE81EFFFFBF77FC008FED1F7F98EFFC00;
defparam prom_inst_14.INIT_RAM_36 = 256'h1B7FFFF9DFFF002FFFDB9FF97FFFC2003AFB398000000E8000062C0080312006;
defparam prom_inst_14.INIT_RAM_37 = 256'h3D3CC00000040000035600002A2001BFFFFFF9087FFFFFFFFDBC3FFFFFFFDFC7;
defparam prom_inst_14.INIT_RAM_38 = 256'hFFFC50BFFFFFFFFF8F13FFFFFFCBAC243FFFFFFFFFC0126AA4EFA99DF708001E;
defparam prom_inst_14.INIT_RAM_39 = 256'hFFFFFFFFF0021BAB3E62E77DC0000E68A1700000000000010A000003C00077FF;
defparam prom_inst_14.INIT_RAM_3A = 256'hB8000002080000B5000002C0001FBFFFFF880FFFFFFFFFF941FFFFFFF3700E25;
defparam prom_inst_14.INIT_RAM_3B = 256'hE46BFFFFFFFFFFA47FFFFFFF2800042FFFFFFFFC00DCBFFE5D18790000078000;
defparam prom_inst_14.INIT_RAM_3C = 256'hFFFFFF00E27A1C424E05E00003F36FCE0000000000006380001B400009FFFFFF;
defparam prom_inst_14.INIT_RAM_3D = 256'h0000400000274000044000005FFFFFC10AFFFFFFFFFFF333FFFFFFE4B41489FF;
defparam prom_inst_14.INIT_RAM_3E = 256'hBFFFFFFFFFFDC5FFFFFFFC802E82BFFFF7FFC00CFF7999109DFC0001E58A9700;
defparam prom_inst_14.INIT_RAM_3F = 256'hFFF0006942070C40C000007BC68B80000000000013E000084000041FFF7FF860;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b1;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'h0000000D900006E0000007BFEFFE1C8FFFFFFFFFFF807FFFFFFF90096107FFFF;
defparam prom_inst_15.INIT_RAM_01 = 256'hFFFFFFFFE0C7FFFFFFE24920C37FFFFFFC0029511006042404007BE6FCE00000;
defparam prom_inst_15.INIT_RAM_02 = 256'h0006904828000000001D7F55700000000000074C0005100000007EFFFE0A07FF;
defparam prom_inst_15.INIT_RAM_03 = 256'h00030600003800000001EFFFC0C1FFFFFFFFFFFD64FFFFFFFC4A03C1DFFFFFFF;
defparam prom_inst_15.INIT_RAM_04 = 256'hFFFFFF1C9FFFFFFF8802F137FFFFFFC080E81004000000001ECD509C00000000;
defparam prom_inst_15.INIT_RAM_05 = 256'hBD0003000260000FBC4DCE000000000001FF00011C000000001BFFE07B3FFFFF;
defparam prom_inst_15.INIT_RAM_06 = 256'h4FC000EB0000000084FFD0323FFFFFFFFFFFEDD7FFFFFFF90502007FFFFFF005;
defparam prom_inst_15.INIT_RAM_07 = 256'hFFF951FFFFFFFF22824847FFFFFC000000010000000003A627D7C00000000000;
defparam prom_inst_15.INIT_RAM_08 = 256'h000000000007C60109C000000000002260005E800000000007840583FFFFFFFF;
defparam prom_inst_15.INIT_RAM_09 = 256'h003160000000080BCD21603FFFFFFFFFFF9C3FFFFFFFE0830884FFFFFF000401;
defparam prom_inst_15.INIT_RAM_0A = 256'hEFA7FFFFFFF80020201FFFFFC00090000000000003EAE40CF000000000001F20;
defparam prom_inst_15.INIT_RAM_0B = 256'h00000003F0D47D7C00000000000E90001B700000000003FBC07A0FFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0C = 256'h2C0000000000FEF00DFFFFFFFFFFFFF871FFFFFFFF8000E05BFFFFF002110800;
defparam prom_inst_15.INIT_RAM_0D = 256'hFFFFFFFFE00002037FFFFC0005300000000003F977889F0000000000079C000D;
defparam prom_inst_15.INIT_RAM_0E = 256'h0001F8FD00CF8000000000033E0006E6000000000045D902607FFFFFFFFFFF64;
defparam prom_inst_15.INIT_RAM_0F = 256'h00000000007C405C7FFFFFFFFFFFE4EFFFFFFFFE4009003FFFFF003080580000;
defparam prom_inst_15.INIT_RAM_10 = 256'hFFFFFFD0201108FFFFC000402000000001E02F93D3C00000000001F180039B80;
defparam prom_inst_15.INIT_RAM_11 = 256'hC0F532E9F0000000000078C001C6C000000000041C401FC3FFFFFFFFFFF02DFF;
defparam prom_inst_15.INIT_RAM_12 = 256'h00000000C602797FFFFFFFFFF8C27FFFFFFFF10002065FFFF000009140000001;
defparam prom_inst_15.INIT_RAM_13 = 256'hFFFE60150A33FFFC0018804000000183F2F08C7C000000000033F000E4700000;
defparam prom_inst_15.INIT_RAM_14 = 256'h8F2D3F00000000001C1800725C0000080000003140BE3FFFFFFFFFFE209FFFFF;
defparam prom_inst_15.INIT_RAM_15 = 256'h000004F009FBFFFFFFFFFF91AFFFFFFFFFEC1806027FFF00030010000005BF4F;
defparam prom_inst_15.INIT_RAM_16 = 256'hF8E40380FFFFC01008000000078FFBFF0CC7800000000006CC001E6E00000000;
defparam prom_inst_15.INIT_RAM_17 = 256'hB3E000000000010F000E370000000000000108C0FF5FFFFFFFFFC937FFFFFFFF;
defparam prom_inst_15.INIT_RAM_18 = 256'h0001344EDBFFFFFFFFF343FFFFFFFFFF2004B085FFF000000000000607AE5108;
defparam prom_inst_15.INIT_RAM_19 = 256'h8D4120BFFC00110800000502C6ED8738F80000000000D1C00713C00000000000;
defparam prom_inst_15.INIT_RAM_1A = 256'h000000000072C001F2A000000000000000F40BD1FFFFFFFFFD017FFFFFFFFFC4;
defparam prom_inst_15.INIT_RAM_1B = 256'h07608B8FFFFFFFF8073FFFFFFFFFFC1200C053FF0000000000027807F624361F;
defparam prom_inst_15.INIT_RAM_1C = 256'h10127FC0040078000060738E5EE5C3E00000000034B001E97800000000000000;
defparam prom_inst_15.INIT_RAM_1D = 256'h0000000EDC00FD1E0000000000000001C41C37FFFFFFFC4D4FFFFFFFFFFF0600;
defparam prom_inst_15.INIT_RAM_1E = 256'h0734DFFFFFF0E02BFFFFFFFFFFA1C080301FF00004000000C03BDC351F98F800;
defparam prom_inst_15.INIT_RAM_1F = 256'h03FC0000000000D00FE3D780E63F00000000075E0039AE800000000000000010;
defparam prom_inst_15.INIT_RAM_20 = 256'h0003E3001EE3A0000000000000000000D9FD7FFFB1FE84FFFFFFFFFFF0080024;
defparam prom_inst_15.INIT_RAM_21 = 256'h07BE4C8573227FFFFFFFF7FD01000A0C7F00000000006023E9E7201EC7E00000;
defparam prom_inst_15.INIT_RAM_22 = 256'hC0000020003A11E098700599F000000000DBC00F25F00000000000000000001E;
defparam prom_inst_15.INIT_RAM_23 = 256'h396007967C000000000000000000016C77DC7DFE783FFFFFFFFBE782E00A0433;
defparam prom_inst_15.INIT_RAM_24 = 256'h77FFE7F40FFFFFFFFF39E0141A30A1F0000010001E847BEC1C00CA7C00000000;
defparam prom_inst_15.INIT_RAM_25 = 256'h0000000628507E730036CF000000001BF801EE9C000000000000000000006422;
defparam prom_inst_15.INIT_RAM_26 = 256'h00F94FC00000000000000000094744E25E7DB98BFFFFFFFEB67802800F06DC00;
defparam prom_inst_15.INIT_RAM_27 = 256'h78FB01FFFFFBFFFBEC29500CC4890000000003AA787FFE800053C0000000066C;
defparam prom_inst_15.INIT_RAM_28 = 256'h0001E63C3F89D86204E8000000012F007E83E00000000000000908D005EAEC80;
defparam prom_inst_15.INIT_RAM_29 = 256'h49F80000000000002FBFFB75C70AE00A67007FFFBF7FEEF2C22E1701E0000000;
defparam prom_inst_15.INIT_RAM_2A = 256'h00DFFFFFEEA61C0001400680C000000000F9EFDFFAAC00813E00000000C9807F;
defparam prom_inst_15.INIT_RAM_2B = 256'h7C7FBBF57B023ACF800000003AE00F8A7C0000000000001FFFA4BFBF7F0F1B7C;
defparam prom_inst_15.INIT_RAM_2C = 256'h801000000001FFFE049FF3EAFE00F80017FFBFF7987000108800200800000000;
defparam prom_inst_15.INIT_RAM_2D = 256'hFFFDFEC394042015014C02000400000FB7EA7FE4000E13E00000000D340FEF3F;
defparam prom_inst_15.INIT_RAM_2E = 256'hFA3E0980D7C4FC00000002EC03F347E80080000000FFFA1C9FFED64DFF000000;
defparam prom_inst_15.INIT_RAM_2F = 256'h20000025FFFC1CAFFFF47B180000001EFE300081A10002A47000000000000754;
defparam prom_inst_15.INIT_RAM_30 = 256'hCC00010020005C40000000000003935F8164603C2C7F00000001CF1BFC33FE40;
defparam prom_inst_15.INIT_RAM_31 = 256'h2BC01E5C9F20000000F5897F4CFF80000000097FFC1BF4FFFEDFA4000000036F;
defparam prom_inst_15.INIT_RAM_32 = 256'h003C7FFC1EC6FFFBC9DD0000000037C08000000000098000100000000383FFF4;
defparam prom_inst_15.INIT_RAM_33 = 256'h000000000170000400000000E6A7FF4E880F01A7F00000001662FFDE3FE10040;
defparam prom_inst_15.INIT_RAM_34 = 256'h0BC113FE000000249B3FE29FFC01000001FFFC0CCAC4E9F0C9F80000001629C0;
defparam prom_inst_15.INIT_RAM_35 = 256'hFFFE0E79117CBF3CF800000000602040000800009B0002800000058FC1CFC82C;
defparam prom_inst_15.INIT_RAM_36 = 256'h000008030000C0000001C78C87D2D501F1DDFF000000035FFFFDE7FF00000009;
defparam prom_inst_15.INIT_RAM_37 = 256'hBA7FC0000003C3FFFE7BFFF00000007FFF07338C94CFE2878000000038800010;
defparam prom_inst_15.INIT_RAM_38 = 256'h8191ABEB41FCE6F00000000C000C000000002051046000000053F289211002A8;
defparam prom_inst_15.INIT_RAM_39 = 256'h00400417B8000000E7ED8008A301785D1FF000000052FFFF863FF400006147FF;
defparam prom_inst_15.INIT_RAM_3A = 256'hF84000003A3F7FE53FEE0000082FFFE1CC10E0070FCE4E000000018400000000;
defparam prom_inst_15.INIT_RAM_3B = 256'h58F90410B995F0000000000000000000000064E0000000EFDE6E200080551E8F;
defparam prom_inst_15.INIT_RAM_3C = 256'h0000E00000002B2F2F201F00083F47FE0000007F2FFFF247FBC4001045FFE0E6;
defparam prom_inst_15.INIT_RAM_3D = 256'h00085F4BFFFED9FEF0480471FFF073E43F82D237A90E00000001000000000000;
defparam prom_inst_15.INIT_RAM_3E = 256'hC5E603713780000000000000000000000000020000222EF2E106A0000BA1FF80;
defparam prom_inst_15.INIT_RAM_3F = 256'h000000001A003D1E05400149D0FFFC000001CDFFFF3CFFFDC0127FFFF8794C7F;

pROM prom_inst_16 (
    .DO({prom_inst_16_dout_w[30:0],prom_inst_16_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_16.READ_MODE = 1'b1;
defparam prom_inst_16.BIT_WIDTH = 1;
defparam prom_inst_16.RESET_MODE = "SYNC";
defparam prom_inst_16.INIT_RAM_00 = 256'h251388F167EBE643CA078A715F23A06F78338494F3EF3E3F80CCD4FFE1F99B79;
defparam prom_inst_16.INIT_RAM_01 = 256'hAE28CC0FE243B0C0F3F367F87E7CF6D975C6583786D2AC900B7325B6A8AC001C;
defparam prom_inst_16.INIT_RAM_02 = 256'h0F5AB76D4F675435AF5D4F2A2B7800F1B96AF39039F472728E811B7F6800E3AB;
defparam prom_inst_16.INIT_RAM_03 = 256'h0F03C369E41CB70283A9AFC07592ECDB1E4574897CC0160CFAE00FF91FD8C509;
defparam prom_inst_16.INIT_RAM_04 = 256'h9E5137BFCF05523D5E3DE641EB0D7DBCB8CB21165C4A71090E699D3ADC1FE00D;
defparam prom_inst_16.INIT_RAM_05 = 256'h0D52D9F36E7558A84B97830F16A6037840B0497A318C47C6EF9E322CA4C5C6AA;
defparam prom_inst_16.INIT_RAM_06 = 256'h1CAE38F85BB81C74D5148FBCB29A2F4E7AC99DE6BC1FF7C74A8068E5759B459D;
defparam prom_inst_16.INIT_RAM_07 = 256'hD9DCE6E189BC262560001AC9FCBE7AD359B019731E0A56F4CDC58986B2996502;
defparam prom_inst_16.INIT_RAM_08 = 256'h4DBC9E90E435A6A0B4187F7DF52A43A97B558A090803A4CA40FED5D2B9EE0B5C;
defparam prom_inst_16.INIT_RAM_09 = 256'hA56142C40169B561B027166C05000821AE4AB7A5800949386062D20D2F59C275;
defparam prom_inst_16.INIT_RAM_0A = 256'h124B1D40071639788DAA24373900145B1E3D30CB88EC9C2E0A1FA77D33732A02;
defparam prom_inst_16.INIT_RAM_0B = 256'hC7C4EE9C426FF380686DEA7BFAC9B555DA309C180E43B611C67CF3DB62E20EC4;
defparam prom_inst_16.INIT_RAM_0C = 256'h8F2745A9B10F7E5058449EA3828BFC8757F6D07EFFB0875EB19303F83B845836;
defparam prom_inst_16.INIT_RAM_0D = 256'h0E89FFBFE283B7FF7AA6B21EC4D64E2194BD20A1CF0A60636068E05BE3BA3E06;
defparam prom_inst_16.INIT_RAM_0E = 256'h45F9252F5EC5513801857777120C61A2047761F5C46C481ED706313EFBC10EEA;
defparam prom_inst_16.INIT_RAM_0F = 256'h37BDE7CAD999B1D114AA62BC2F45E1E26ECB54871D27F48731C2D2C02C301F24;
defparam prom_inst_16.INIT_RAM_10 = 256'h7D057E39533B6E4E1886B97D423A03F749C45CC86D7CD550EA078528199C7ED9;
defparam prom_inst_16.INIT_RAM_11 = 256'hE1F038ABA02B0E41047EE1F9D72FB6746F16E56AC89779C7069B2B3894B52427;
defparam prom_inst_16.INIT_RAM_12 = 256'hB73FB44EA684884F0C9C1E5658D19C07A1FFA570603EEB0B75A2F6F29B3A8E42;
defparam prom_inst_16.INIT_RAM_13 = 256'h7EF28E80113C8F0D7C94406AB7F2D09FEA25DC41B81ABF820EF31982B908CE3F;
defparam prom_inst_16.INIT_RAM_14 = 256'h5C6C9E5B865D8EE1958DB2351817AB8DC92E06C3567CF62242B7918939E43EAE;
defparam prom_inst_16.INIT_RAM_15 = 256'h2BB3DBCD6F8C0288D330E7617998029D68E3A6206E130F4B9CE4240FFE25FC7D;
defparam prom_inst_16.INIT_RAM_16 = 256'hA683326AB212FFE84A3947678477131913271A81CEBCA9C3AC88C64509EAFAE2;
defparam prom_inst_16.INIT_RAM_17 = 256'h6BA821057F59F51C5DC5318ABC5069D4C73AC5279DCDDE969292D0EF6B9D01FB;
defparam prom_inst_16.INIT_RAM_18 = 256'h2DBA94396EE9029358E1E3A43C4EF2A271C0D7D9BD889050D8383AB4094EE769;
defparam prom_inst_16.INIT_RAM_19 = 256'hE7D379A48503250AA9A644A671094FEA3F048D7DF8B8F5D0073BAE23E7B91558;
defparam prom_inst_16.INIT_RAM_1A = 256'hF58CE0E5FB354AFA2D181050F6795854D2DE2825B69B0352244D8DBC0072A084;
defparam prom_inst_16.INIT_RAM_1B = 256'hD7B60B214ABF43E1EBAC5F98638EC60F91FB889C839176770BE496866F59F547;
defparam prom_inst_16.INIT_RAM_1C = 256'h0F6AD94569EC22AF7E661091E13B6BF97FF547C63BBB805238F503189A42AF37;
defparam prom_inst_16.INIT_RAM_1D = 256'h028A0B434F946BDD3F00D1A994B768D71E28BE3C8D865338F90F4DF8454945FE;
defparam prom_inst_16.INIT_RAM_1E = 256'hDF4BBCBE51CA01601ED3404DA90F600C43BFE0557B2F0C21FE12DF3D7D092D3E;
defparam prom_inst_16.INIT_RAM_1F = 256'hA71505B3180A7E97DA8980E241F0F58424C51DA4721E4600BF4A1AA20C3F8900;
defparam prom_inst_16.INIT_RAM_20 = 256'h4A0AC396E38EC0A4C7A3AB816EDFF7F0CC6B8231CEAA7B4BD4F5F5452130522A;
defparam prom_inst_16.INIT_RAM_21 = 256'h083EBFBA12173FF4A57F90C8CFFCF2D5F361413377A45099341A9E58B7CC7FC4;
defparam prom_inst_16.INIT_RAM_22 = 256'h9018F7137C33A928DE6CFAA1F01FF0306C99FADFE893F30B80ECE7E1832C72E2;
defparam prom_inst_16.INIT_RAM_23 = 256'hD920CA981D49A3EA783EA5CED3BA386E1EF81A7FE36CF4450F040EA848DA8DDD;
defparam prom_inst_16.INIT_RAM_24 = 256'h905E1121142E58C9DD87C3943AE6EB1C112BA9A65318B5295F26C8D2354F8334;
defparam prom_inst_16.INIT_RAM_25 = 256'hF8C99BC80F0CA488416604051FC3E297801466530F169B1C0B2DE12BB711A65C;
defparam prom_inst_16.INIT_RAM_26 = 256'h3976909BC3DD9E87AB21537E1ED61B81F809D283A67A9C9F08E170179676BA83;
defparam prom_inst_16.INIT_RAM_27 = 256'hAF795A789A7C19AF67972780C297B22B2CCE49B156BD568E568414BE5726B5AE;
defparam prom_inst_16.INIT_RAM_28 = 256'h1EAE4A433E683880FC03A1C06908A09C94C4F07FBF2276A0C84D194520BA88D1;
defparam prom_inst_16.INIT_RAM_29 = 256'h8E003BFA468799617172B87E4A9F2398BB6CDE2BC3244E4784C003FE1720DBFD;
defparam prom_inst_16.INIT_RAM_2A = 256'h7FE62893ED9CF6F82A0944D94CD67CB4E098743A20BEACCDB17F89F8A40F2B3E;
defparam prom_inst_16.INIT_RAM_2B = 256'h2C6256CE9FAA9D3D8B0195F383A4243AC53B03FEC0B90385E3DA532B29634028;
defparam prom_inst_16.INIT_RAM_2C = 256'hC7F8F3211E34EF272905198517D609E6F2E3E79A0CB9F833D736C53FD40C4ECE;
defparam prom_inst_16.INIT_RAM_2D = 256'h5DCC61C8B05C2C005F062B1D3F3AB3B1E73A4F0A8C4D9CC11EB2C6CD7F26622B;
defparam prom_inst_16.INIT_RAM_2E = 256'hFC78B043A0D003473D2F261C311CB5E02E7939BDB362570A3D9E436F0E5B3887;
defparam prom_inst_16.INIT_RAM_2F = 256'h9730DC7B601DD2E5AAC5D7AFCFDC3E67A6CFDFBD37F5F50EB948283AD59AB3D2;
defparam prom_inst_16.INIT_RAM_30 = 256'hBAEFC3DE0BEA54D6D4442A8A273CAA1F3F1AAA44A3465383BD43AC545E6AAEC1;
defparam prom_inst_16.INIT_RAM_31 = 256'h72A9F16C2F8EF0C33FF2D1FA2907E61FAD573008D432EBCF06FD77A6080E6EA6;
defparam prom_inst_16.INIT_RAM_32 = 256'h409F44DB98D3C4380D1CC5CDFC06E21D0DB837C3A92055BCCBF44AEC8F7BE3E4;
defparam prom_inst_16.INIT_RAM_33 = 256'hE468177F590E5CA58C7FEA1C4C6848F723EFC313EE60132E005C797BA9F5BFDB;
defparam prom_inst_16.INIT_RAM_34 = 256'h90F226F91D25511ECEA1E1B029DF7F5A78F0255A7AB734781B6CBA8B645568C1;
defparam prom_inst_16.INIT_RAM_35 = 256'h5A48E65D13D48E625D8CF10435839F0553DDE04FD21751A9CF68518EEABC9903;
defparam prom_inst_16.INIT_RAM_36 = 256'h4504CB13F66678AF8B5A0DEFF97648345BF7BF0777D7EDEBD890FE068FF7FF06;
defparam prom_inst_16.INIT_RAM_37 = 256'h7AC90CCEB672B530D4578463945CF040040DA7D18719E20F11E9D3B9A98C2D17;
defparam prom_inst_16.INIT_RAM_38 = 256'h4392C99380A7C13976A4EE776A50B09F90B2013779E70B0DDFE3D667B0FA4A73;
defparam prom_inst_16.INIT_RAM_39 = 256'hA91075A9017CCFB25F0D02698B5ACC44E40C8A2FBB8807E8996228EE019618B1;
defparam prom_inst_16.INIT_RAM_3A = 256'h1E23D250FE8A05E8A855341847E2B664E46A3D5766BB498ADFBAC2863295C908;
defparam prom_inst_16.INIT_RAM_3B = 256'hB64DF0D2EBFC34B46F5BA78BBDD5BFCB3FB185C92334D84962CFE6D82453F204;
defparam prom_inst_16.INIT_RAM_3C = 256'h1BAAB54A1560B1F6FE0A6250388A23E3AB59B06CA90572C863B047856593AC8A;
defparam prom_inst_16.INIT_RAM_3D = 256'hFAF6535E49E0D8A157C7944DE76B8EC2645A9CF2419E63EB19B2D74A968A27AB;
defparam prom_inst_16.INIT_RAM_3E = 256'h9A5E0338AABB05C34BEECBD0A0F6FAF19EEE3A7944980B731A0CBC0C7F4BCED9;
defparam prom_inst_16.INIT_RAM_3F = 256'h3EFB4E29C83D85381C92E8E45F43B127F97491570F5E17594D8D9AF6FB834C46;

pROM prom_inst_17 (
    .DO({prom_inst_17_dout_w[30:0],prom_inst_17_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_17.READ_MODE = 1'b1;
defparam prom_inst_17.BIT_WIDTH = 1;
defparam prom_inst_17.RESET_MODE = "SYNC";
defparam prom_inst_17.INIT_RAM_00 = 256'h01D7860194EA1743CA3DFC621B36684D53DCD72A7810FC007FF32A4006040C80;
defparam prom_inst_17.INIT_RAM_01 = 256'hEFACB2F49DBF800F0C0C10000101082C81D5EF2665B442077DB43216A9780104;
defparam prom_inst_17.INIT_RAM_02 = 256'h00A53769F4FB91D61B90C2661F7C00F1CF8903F0EB8BB2F2FDFC1DA9D3B06260;
defparam prom_inst_17.INIT_RAM_03 = 256'h4503F41E61FFF3E77C2ED4A7838558DEDFDBC6B0832801F20000000000270800;
defparam prom_inst_17.INIT_RAM_04 = 256'hBDAE958037002D8042580000087100B84F0F0C15E1BF985AE497D343DC01C076;
defparam prom_inst_17.INIT_RAM_05 = 256'h4EA9846DEF627B8BFC1C8CFF06E61C79403DD9994FACFFFD142BCF37D0346B8A;
defparam prom_inst_17.INIT_RAM_06 = 256'h1BF66807BFFFEB171C89249C0D13D3F562E382317C0000030000040080000543;
defparam prom_inst_17.INIT_RAM_07 = 256'h6342993D9040A42000001800089E800447F5829D77A03BB10302F998279EBCD8;
defparam prom_inst_17.INIT_RAM_08 = 256'h791B7F0D240ABC738DF7FFBDFF27B7AEA30380FCFFFC070CD6F220C205F2165A;
defparam prom_inst_17.INIT_RAM_09 = 256'h90E0FF7BFE81C65C06C61E010104E4306C45497D8039481860204201275403B7;
defparam prom_inst_17.INIT_RAM_0A = 256'hF81473C00716FB7888886D373C80C052FB83128B823E77E277FFEF7FD936EFC9;
defparam prom_inst_17.INIT_RAM_0B = 256'h1A6F368CE71BE9839E7DFF8D7BBBC57D9A1F6FFFF2F321C1C5D6422343E84EC0;
defparam prom_inst_17.INIT_RAM_0C = 256'h81DEEA51BFCABDD08122B0C123BAD7BD20013836FF32D75EB19353FF03E8742F;
defparam prom_inst_17.INIT_RAM_0D = 256'h0037DF3FFBDBF7DF7AAF3CDEBD39815E700DA004312EE39CBFFF81689F4F131E;
defparam prom_inst_17.INIT_RAM_0E = 256'h1BF90DC6CB300AC7FFB9BFECC3A857A1FBDC91FE76F9D851D778602899B6D74A;
defparam prom_inst_17.INIT_RAM_0F = 256'h980020AB4E8464A873184047D7E6BBE0413BC7F8FB7F7F57BDFB32D9EEF5A7DA;
defparam prom_inst_17.INIT_RAM_10 = 256'h56EE8077FBEFFBED6F7FAC063A0F688979026A945C036EAF5438FB1E3395FD26;
defparam prom_inst_17.INIT_RAM_11 = 256'hB0C33607B194753E1279CC71255F998E801F05381F32EEC0C2704465E95C0C03;
defparam prom_inst_17.INIT_RAM_12 = 256'h07C3227E0388CB136B778E048FA5CC0014003AFFDFFFFB8F80AB614E66658366;
defparam prom_inst_17.INIT_RAM_13 = 256'h8011777FE66F7AF1BB5893C139873E000631F5C040E5408C3C101C3447002180;
defparam prom_inst_17.INIT_RAM_14 = 256'hD7AE7E1111A00B422C06AB90F820400FF14AE2839839F5CC7CFF413380A30CA8;
defparam prom_inst_17.INIT_RAM_15 = 256'h32C909B682BAC0DE92AD56578767F012806459DFF1EDB04FE314E0F481CF801C;
defparam prom_inst_17.INIT_RAM_16 = 256'h665FED9D0D42E3F01838B8B07BE80BFB1D9F0802003F21C9AD347E3F001083FC;
defparam prom_inst_17.INIT_RAM_17 = 256'hA79801005FED56DD914B0F8840007E18A89C90769399DF1CBCB404AD8F601004;
defparam prom_inst_17.INIT_RAM_18 = 256'hCFDEC15FA1E78780CA2AF0E103C6C802261A28241988DE61A403C54BFE109D46;
defparam prom_inst_17.INIT_RAM_19 = 256'h18298008053ED9710679BB5FAF5B8479FF04811FD184BFE20AB9ECA001BE8EAF;
defparam prom_inst_17.INIT_RAM_1A = 256'hF58CE5F9B4ADF1757CF800117F81ADF9DED15E4F18C8157457C418D8FFF21104;
defparam prom_inst_17.INIT_RAM_1B = 256'hD03398FCB7C30FFCBD40230FDF8243008A0C009CF5E2242ABE67FF75E7D244FF;
defparam prom_inst_17.INIT_RAM_1C = 256'h984882DF989140FFBFF417B81F4556FCFFF7F8ED65FC9ECADEF5035960736BD7;
defparam prom_inst_17.INIT_RAM_1D = 256'hBFF508FD733C4787BF00D1D41AD01B70CC5B7879B74B06D792B68D23C4584420;
defparam prom_inst_17.INIT_RAM_1E = 256'hA8FB9564EC771CCAC2A28DBD880F400013A7E5E2E4135920FE13D4E29D962D7F;
defparam prom_inst_17.INIT_RAM_1F = 256'hB758761C41C6741FDAA52E47A237FDEFFB07469B3565C3FFB75BE50791CC6C8F;
defparam prom_inst_17.INIT_RAM_20 = 256'h037F64151C683FFDCFBC41E7D2E29DB40F1B4E04BA6168B25C3943C16170522A;
defparam prom_inst_17.INIT_RAM_21 = 256'h67F24C4FD751AEC80F4079C85EDC625DFF5F925EFEB0001B888642294FFFFFBB;
defparam prom_inst_17.INIT_RAM_22 = 256'h77E0CA3B63B461193EDCEE1FFFFFEFC3B4E81E679C2CCF7FFF10F949B92C9412;
defparam prom_inst_17.INIT_RAM_23 = 256'h4303682702BE7FF5801D200C52B85513DD2F247A74CA7774221BEFAB58D83FD5;
defparam prom_inst_17.INIT_RAM_24 = 256'h2C400DEA06DA8D32806EA7F63AF8EF3FED3272D5B0C2048ABB85C7FBCAF003DE;
defparam prom_inst_17.INIT_RAM_25 = 256'h3B43E93CA3AD03B9A2E1FFFAE003954043C629D0F0FDFDC00AC96010956E5C76;
defparam prom_inst_17.INIT_RAM_26 = 256'hD7F370601CA26007F2259ACFA510A13F0B8F204AE265A01F377FFF77FE7FF46C;
defparam prom_inst_17.INIT_RAM_27 = 256'h0B2FB9F1176A6B8099F4B7FFFFFAC5C38DA23FF246CA1317307BEB0007537E56;
defparam prom_inst_17.INIT_RAM_28 = 256'hAC017849EC20A3100BFC00009076B3EE519C0F0040F4003CE9D68707EE8D1A9E;
defparam prom_inst_17.INIT_RAM_29 = 256'hC380100439039E85CDEA761A8EFFFC8A754DB371C3093C22FFB7F9FEB8CF20F0;
defparam prom_inst_17.INIT_RAM_2A = 256'h69E408ECE41FF057D9FFFBA0B1207F27333045D39AA2A4024E0009C10B92D2C5;
defparam prom_inst_17.INIT_RAM_2B = 256'hA0451A6F9A2782C03203E98F6181AED9C0020000403FFA2B898E453F5544F611;
defparam prom_inst_17.INIT_RAM_2C = 256'h870180051FF8CB5FFFA8A87DFB95A380ACAE75333FF0868D3ECD1AA0080F8C92;
defparam prom_inst_17.INIT_RAM_2D = 256'h9E11E60E5423C31FA0F210891BC2C665F38DD5B5DD4080081FACECD75FF7A67B;
defparam prom_inst_17.INIT_RAM_2E = 256'h71BF4B98E04001476A344D9DD65D8DF0024039FDBC6C8772E17AFE12DE8CF23E;
defparam prom_inst_17.INIT_RAM_2F = 256'h0611FCFF8386B341AA886F1593124129EF9721CBE4021A998014080AFA14A6C9;
defparam prom_inst_17.INIT_RAM_30 = 256'h06D9F03E404A2028000420BFC7891647A2CF2675A34457E4302DA5937727FEC0;
defparam prom_inst_17.INIT_RAM_31 = 256'h13A73D446F8FDF0C7CC61BAE5AEFE61FAD7FFFF0E759E75231E67D6E732FC22F;
defparam prom_inst_17.INIT_RAM_32 = 256'h5FF7FA9CED5AF4A6693CAB4754B0F34E54657BC161C0B00CC2FD5F80B592B819;
defparam prom_inst_17.INIT_RAM_33 = 256'h5398D670790E1E26FC37D59F0EB231DD6F1FC313EFFF8004436D96F67FF5BFDB;
defparam prom_inst_17.INIT_RAM_34 = 256'hBFF237FBF6959AE1EBAF848BEDDF7FFBBFFF468CB6A4C0837C58B781FDE983C0;
defparam prom_inst_17.INIT_RAM_35 = 256'hFDB0F090627EDFC21FCB32FC3281379001BFF84FD2154DE95ED7A1F0AC60B08F;
defparam prom_inst_17.INIT_RAM_36 = 256'h1BF54332F79B7FFBE9A00F2E768FA40B5BFFFF7BC8E5648ABB9131FBF7FBBCFF;
defparam prom_inst_17.INIT_RAM_37 = 256'hFEFEDF303A5E102F33507FBFDFBF1FFFB80E3B282202BF0072EA330B3F447477;
defparam prom_inst_17.INIT_RAM_38 = 256'h2B4332CD93B1E3857D4536F286AE24EE77FAE99777EEFEF320C1FA78001E33F7;
defparam prom_inst_17.INIT_RAM_39 = 256'hFF67FC7FFE9FF004130B806F470DFCFFEBE3614CD5A6691E361D7FFFFE79E74E;
defparam prom_inst_17.INIT_RAM_3A = 256'hD098039ACB72AF66A7AEFBE7981D4986E873ACCAF94777A12A364C77B7D41D9F;
defparam prom_inst_17.INIT_RAM_3B = 256'h07004282FA3E3790EA4909E97B98A0E9F0BFFF36CBFF0C0141F806E819FFFFFF;
defparam prom_inst_17.INIT_RAM_3C = 256'hE675CBB0EA50B9E2FBB4022BDDFFDC18100183D59C12D2C41D5FB87A026C000F;
defparam prom_inst_17.INIT_RAM_3D = 256'h12F9633F8E72F840E0080B8018060FFC789C1FF639AF9DFDBBDEFC1BA738DC74;
defparam prom_inst_17.INIT_RAM_3E = 256'h1C89D04787AFB20EF069D3EBE109859FE518C454140C0A7FF57002FBF3940100;
defparam prom_inst_17.INIT_RAM_3F = 256'hC1001189C92187FBE3651F1BA0100001FF877165FFCE4800200000000000FF97;

pROM prom_inst_18 (
    .DO({prom_inst_18_dout_w[30:0],prom_inst_18_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_18.READ_MODE = 1'b1;
defparam prom_inst_18.BIT_WIDTH = 1;
defparam prom_inst_18.RESET_MODE = "SYNC";
defparam prom_inst_18.INIT_RAM_00 = 256'h01F3BFFE3565F743CA3FFF8392ED276A03DB39F6D80003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_01 = 256'h6FF4FE7280007FFFFFFFFFFFFFFFFFF7FE00003CFE947091FA9E18E5A7F80004;
defparam prom_inst_18.INIT_RAM_02 = 256'hF000306F4FCFD17BE81592E1FF7800F1F7C7FC1D587FF2F2FFFFE1CD54DB9361;
defparam prom_inst_18.INIT_RAM_03 = 256'h34FC07161FFFF3E7FFD0E6F61A7960FEA5EAEE300017FFFFFFFFFFFFFFFFF7FF;
defparam prom_inst_18.INIT_RAM_04 = 256'h20D48B8000FFFFFFBDE7FFFFF7FEFF44000CBDC7FC7F681A0D28B0FBDC01C079;
defparam prom_inst_18.INIT_RAM_05 = 256'h0F97E47FC70E450355CC7FFF06E61E213FC11387FFACFFFFE0332A2EFE304B9B;
defparam prom_inst_18.INIT_RAM_06 = 256'hE0C4E7FFFFFFFFE818D5E7FFD01BDFDF89F7F80003FFFFFCFFFFFFFFFFFFFA00;
defparam prom_inst_18.INIT_RAM_07 = 256'h9D4280026FFFDBDFFFFFE7FFF7614007BA55EBF4BE224B96973FFD98279F2647;
defparam prom_inst_18.INIT_RAM_08 = 256'hC9089E4064079DA183FFFFFDFFCF105037B07FFDFFFFF80F62D17DE409F01DA8;
defparam prom_inst_18.INIT_RAM_09 = 256'hAC1FFFFFFFFE07969FC31E010706E106DF4000027FC6B7E79FDFBDFED8A003DE;
defparam prom_inst_18.INIT_RAM_0A = 256'h6E00003FF8E944877777D2C8C000E2AE00811EE38070E161FFFFFF7FE30E100F;
defparam prom_inst_18.INIT_RAM_0B = 256'h006EDE8C0DBC587FFE7DFFF1BD8406DB85FFFFFFFD03C55FCCF6420343A81229;
defparam prom_inst_18.INIT_RAM_0C = 256'h7FFFFFFE41F3652F158240A163FDF368600007C900CD28A14E6CAC0003F24C03;
defparam prom_inst_18.INIT_RAM_0D = 256'h00002040042408008550421EFA57B1C00005A0135DC61FFFFFFFFE45600FBA81;
defparam prom_inst_18.INIT_RAM_0E = 256'h39F90215710FFFFFFFFE325C03EF305FFFFFFE0078A6CDA9A7702008D9D29962;
defparam prom_inst_18.INIT_RAM_0F = 256'hFFFFD8AC6861DF595010043057755F604004380000808028420402DE51F67000;
defparam prom_inst_18.INIT_RAM_10 = 256'h40000000040000100003AF9BFA78000AB9014A2EC3FFFFFFFFCC3700244C03FF;
defparam prom_inst_18.INIT_RAM_11 = 256'hA0332BA04FFFFFFFE31DC07C33007FFFFFE006B26CAFF1C402040B870535EC03;
defparam prom_inst_18.INIT_RAM_12 = 256'hF803C4E5DF8DF9000201F7EA790D4C00000020000000006000AB86FE03BCC1F4;
defparam prom_inst_18.INIT_RAM_13 = 256'h00110000088000013BE1FFC000011C001CF4EC3FFFFFFF707C701E45C0FFFFFF;
defparam prom_inst_18.INIT_RAM_14 = 256'h966A01EEFFFFF0721C07197007FFFFF00173581BD3AB240043FEFEC48A2F0CA8;
defparam prom_inst_18.INIT_RAM_15 = 256'h3CD5D864027E8000D3ADF8F9A1E3F000006000000000004FFC57E000001E8003;
defparam prom_inst_18.INIT_RAM_16 = 256'h660000000002E3FF90F8000000A0046B3080F7FFFFC02927ADDDDE00FFFF7C00;
defparam prom_inst_18.INIT_RAM_17 = 256'h6067FEFFA00E8DDDE5E70077FFFF801F342EF0A71BE1E030C0B7E0A336FC0000;
defparam prom_inst_18.INIT_RAM_18 = 256'h0DF89300A46838080A74E0BBBFC6C002200000000988DF857C00000000017AFB;
defparam prom_inst_18.INIT_RAM_19 = 256'h00000000053FE1DF0000000000BB6D5800FB7EE001167FFC49B8135FFE400FCD;
defparam prom_inst_18.INIT_RAM_1A = 256'h0A731A01C49DFEB2FC07FFEE8001F1403E9824184709E0881788F547FFF21104;
defparam prom_inst_18.INIT_RAM_1B = 256'hB9705E14C0F8F400B0D263F7FF8243008008009CF7FC5FE0400800001F12AC00;
defparam prom_inst_18.INIT_RAM_1C = 256'h084880DFFF1990000009E84B05EB4003000800F5A7FF23BA010AFCA6007C442B;
defparam prom_inst_18.INIT_RAM_1D = 256'h40000C8AFCD65F8040FF2E001F1A7B7D46020DAD7BCDF844A29022FFC4584420;
defparam prom_inst_18.INIT_RAM_1E = 256'hE8122D5F74F8E1ADC265BFFD880F400003A7E7F7069102DF01EC2CFE90809280;
defparam prom_inst_18.INIT_RAM_1F = 256'hA75977E09D218BE0257D73DF6008021000067A7FC553C00048A40007E2B1AC35;
defparam prom_inst_18.INIT_RAM_20 = 256'h0382DFE255E80002304001F992CE5F1809569DA4FFD47C022EC7BFC16170522A;
defparam prom_inst_18.INIT_RAM_21 = 256'h1EF3440FF898DE826BBFF9C85EDC625DFF7FFC645A7FFFE47D5EED9800000000;
defparam prom_inst_18.INIT_RAM_22 = 256'hFFFF0C952D6FDEF85278660000000003C2A7E0BD7C0000800000FE73BBF1092A;
defparam prom_inst_18.INIT_RAM_23 = 256'h68FC509F00000000001FC6BDA4809EF865FF047F86E9AA9CD1FFEFAB58D8BFDD;
defparam prom_inst_18.INIT_RAM_24 = 256'h7C400DD1248C22DB7FFFE7F63AFEEF3FFEC3B7314E3FF90F1793C004000003E5;
defparam prom_inst_18.INIT_RAM_25 = 256'hC4728B52A52DF3FBE9E000000003F90A3C1CA7D0000000000BF1B7E0DBDFE067;
defparam prom_inst_18.INIT_RAM_26 = 256'h1120F00000000007FC377FF5EAEBB80B880FFCC61594F910FFFFFF77FE7FFFFF;
defparam prom_inst_18.INIT_RAM_27 = 256'h0B3E310BE538547FFFF7B7FFFFFFFFFC0AC59A89A09B6F3AF0000000077D86C1;
defparam prom_inst_18.INIT_RAM_28 = 256'hC9675A8566F0D17000000000FE30100CA47C00000000003F0E8E899237FF9B4A;
defparam prom_inst_18.INIT_RAM_29 = 256'hBF80100000039FF997185A89DEE3F1883E8986FD730C83FFFFF7FBFFBFFFFE01;
defparam prom_inst_18.INIT_RAM_2A = 256'h0A7B7F5965A00FBFFFFFFFFFFFFF8039B6C1F0FA09D39C00000009FE28D60321;
defparam prom_inst_18.INIT_RAM_2B = 256'h6AC42E9B049F80000203FE150C81CD47C0020000403FFC32D920C82B46749003;
defparam prom_inst_18.INIT_RAM_2C = 256'h870080051FFF0C6A644025AFFDB6C3E1FA9F95723A0F7FFEFFFFFFFFFFF00F1B;
defparam prom_inst_18.INIT_RAM_2D = 256'h43E5540D13DFFFFFFFFDFFF7E402FBB458294BC9434080001FBF09D63FC0C1FB;
defparam prom_inst_18.INIT_RAM_2E = 256'h4B1CFD47E04001477FC6E0C5E3147DF0024039FDBF90E1B48F03D6B1E6487CE6;
defparam prom_inst_18.INIT_RAM_2F = 256'h0611FCFFFC18D943F50C2E45571C6506520901381FFFE7F77FFFF7F5001F3B76;
defparam prom_inst_18.INIT_RAM_30 = 256'hA509EE01FFBDFFFFFFFBDF4007F1DB53249561F4A34457EFC1BF73E7551FFEC0;
defparam prom_inst_18.INIT_RAM_31 = 256'h9660FD446F8FFFF05CE7E372C7EFE61FAD7FFFFF079D5F09FC448D70F63349F1;
defparam prom_inst_18.INIT_RAM_32 = 256'h5FFFFF60F196336F9E34EC787C937C4DC03FF03EDE3FFFF33D02A000BA1CCCE0;
defparam prom_inst_18.INIT_RAM_33 = 256'h0458298F86F1E1D90388001FF0C3812CE0FFC313EFFFFC3705313ED1FFF5BFDB;
defparam prom_inst_18.INIT_RAM_34 = 256'h7FF237FBFFFA1C9754FF4C7BEDDF7FFBFFFFF80F3BEB82FB3418E00FB41E3B30;
defparam prom_inst_18.INIT_RAM_35 = 256'hFFFF00E1B60FDF9F178DAC656F498C41A38007B02DEAB216200001FF0F800F80;
defparam prom_inst_18.INIT_RAM_36 = 256'hD00ABCCD0860800014000FD07FFF83FF5BFFFF7FFF06872527930FFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_37 = 256'hFEFFDFFFC29023C9E8CFFFFFDFFFFFFFFFF03C31621FBF03F326C160CD82ED54;
defparam prom_inst_18.INIT_RAM_38 = 256'hFC03C3139E708F7D72EF298B71208E76080516688810000000C1FD800001FBF7;
defparam prom_inst_18.INIT_RAM_39 = 256'h0088028000000000130FFF9030FFFCFFEFFFFFF0E4B5F3F1F1FFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3A = 256'hFFFFFC1C7AFCBCFD5FFFFFFFFFFFFFFB107C313E0E2D67A1753320B650142F80;
defparam prom_inst_18.INIT_RAM_3B = 256'h07F19783844934802AB421AC01AF6014000000000000080141FFF917FDFFFFFF;
defparam prom_inst_18.INIT_RAM_3C = 256'h000000000040B1E2FFFFFDFFFDFFFFFFFFFE439C7FBA463FFFFFFFFFFFFFFFF0;
defparam prom_inst_18.INIT_RAM_3D = 256'hED007CFFE29DC7FFFFFFFFFFFFFDF0007F1C7191CFFF1DE3C798CFF458080000;
defparam prom_inst_18.INIT_RAM_3E = 256'hE0E4D3BCCDAFCDF1E2A6AC033B00008000000000040C0A7FFFFFFFFFFFFFFEFF;
defparam prom_inst_18.INIT_RAM_3F = 256'h00000009C92187FFFFFFFFFFFFFFFFFE0007F17CF341FFFFFFFFFFFFFFFF0017;

pROM prom_inst_19 (
    .DO({prom_inst_19_dout_w[30:0],prom_inst_19_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_19.READ_MODE = 1'b1;
defparam prom_inst_19.BIT_WIDTH = 1;
defparam prom_inst_19.RESET_MODE = "SYNC";
defparam prom_inst_19.INIT_RAM_00 = 256'h01E2FFFFCF1FF743CA3FFFFC1CEA9FB2FF343602180000000000000000000000;
defparam prom_inst_19.INIT_RAM_01 = 256'h9122A1A48000000000000000000000000000003D0295EE80BB9064CC5FF80004;
defparam prom_inst_19.INIT_RAM_02 = 256'h000034904FCAF0E7E00BE61FFF7800F1FB5FFFE1C7FFF2F2FFFFFE0E7927FD1E;
defparam prom_inst_19.INIT_RAM_03 = 256'hA3FFF9F1FFFFF3E7FFFF073A81FEDF014E083DB0000000000000000000000000;
defparam prom_inst_19.INIT_RAM_04 = 256'hC2D6DF80000000000000000000000000000E0207FC8FFCE80A4D8FFBDC01C07E;
defparam prom_inst_19.INIT_RAM_05 = 256'h0F40147FDCA5C6829943FFFF06E61F8CFFFE287FFFACFFFFFFC3C94AFFCFA454;
defparam prom_inst_19.INIT_RAM_06 = 256'hFF0A1FFFFFFFFFFFE0E7917FE7FC20087EDFD800000000000000000000000000;
defparam prom_inst_19.INIT_RAM_07 = 256'hCBBE8000000000000000000000000007DC150BF2512203E730FFFD98279FCD3F;
defparam prom_inst_19.INIT_RAM_08 = 256'h4949FE242407A1C87FFFFFFDFFF7CFFFC48FFFFDFFFFFFF07BC47DF3F60DE141;
defparam prom_inst_19.INIT_RAM_09 = 256'hE3FFFFFFFFFFF818ECC31FFEFBF90E93D8C000000000000000000000000003EB;
defparam prom_inst_19.INIT_RAM_0A = 256'hCE00000000000000000000000000FDE2040105D3817BFB1FFFFFFF7FFD31FFF2;
defparam prom_inst_19.INIT_RAM_0B = 256'h4076EE8C6EFEC7FFFE7DFFFE7C7FF8087FFFFFFFFFFC06781AB63D7CBC17EB3E;
defparam prom_inst_19.INIT_RAM_0C = 256'hFFFFFFFFFE03B727E1FD7F5EFC4E607DE0000000000000000000000003FDFC20;
defparam prom_inst_19.INIT_RAM_0D = 256'h00000000000000000000001EFF5F8020010DA00FADA1FFFFFFFFFF951FF0067F;
defparam prom_inst_19.INIT_RAM_0E = 256'h09F901EB68FFFFFFFFFFC143FC010FFFFFFFFFFF80C927FE988FEFD726A9E23A;
defparam prom_inst_19.INIT_RAM_0F = 256'hFFFFFF5072ACFFFCA7EFFBDFB8D92A604000000000000000000002DFA7F21000;
defparam prom_inst_19.INIT_RAM_10 = 256'h40000000000000000003AFE5FA2800039900310A3FFFFFFFFFF190FFC343FFFF;
defparam prom_inst_19.INIT_RAM_11 = 256'hA00D629FFFFFFFFFFC343F8190FFFFFFFFFFF83CD7FFF7BFFDFDF7FBF9D4AC03;
defparam prom_inst_19.INIT_RAM_12 = 256'hFFFC07599F8F75FEFDFBFFFFB548CC00000020000000000000ABFB7E013C4000;
defparam prom_inst_19.INIT_RAM_13 = 256'h00110000000000013BFE1FC0000020000362A3FFFFFFFFFFBE0FE0CC3FFFFFFF;
defparam prom_inst_19.INIT_RAM_14 = 256'h0BB9FFFFFFFFFF8A83F8230FFFFFFFFFFE8396C7D293AAFFBDFEFFF8173F0CA8;
defparam prom_inst_19.INIT_RAM_15 = 256'hC0E4C5E4C33C3FDF53EDFF9FF6EFF000006000000000004FFFBFE00000008000;
defparam prom_inst_19.INIT_RAM_16 = 256'h660000000002E3FFEAF8000000200008A47FFFFFFFFFD2205210C1FFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_17 = 256'h1FFFFFFFFFF0CC2206A0FFFFFFFFFFE03968D0F713A61FB080B7FD16D8FC0000;
defparam prom_inst_19.INIT_RAM_18 = 256'h591AD4E0A617D0080A7F2A4AFFC6C002200000000988DFF87C0000000000026D;
defparam prom_inst_19.INIT_RAM_19 = 256'h00000000053FFE3F000000000005C1C7FFFFFFFFFE1200019847FFFFFFFFF00E;
defparam prom_inst_19.INIT_RAM_1A = 256'hFFFFFFFE1582008603FFFFFFFFFE019560CFFC0841F0040017F1FF2FFFF21104;
defparam prom_inst_19.INIT_RAM_1B = 256'h198FC106B8040000BE090CFFFF8243008008009CF7FF9FE000000000006F23FF;
defparam prom_inst_19.INIT_RAM_1C = 256'h084880DFFFE2F00000000007D378BFFFFFFFFF0360003D85FFFFFFFFFF80754C;
defparam prom_inst_19.INIT_RAM_1D = 256'hFFFFF1980012C07FFFFFFFFFE01CD38AC9FE9C32003000470230AFFFC4584420;
defparam prom_inst_19.INIT_RAM_1E = 256'h17F5C2C04B0001D2C2EC7FFD880F400003A7E7F7F8AF0000000002A1647FFFFF;
defparam prom_inst_19.INIT_RAM_1F = 256'hA75977FF1CE0000000039A051FFFFFFFFFF8660006F03FFFFFFFFFF8032AF33C;
defparam prom_inst_19.INIT_RAM_20 = 256'hFC29C003AC17FFFFFFFFFE01E79F050FF71A385B000073820BAFFFC16170522A;
defparam prom_inst_19.INIT_RAM_21 = 256'hFEB3A3F0001F61013BFFF9C85EDC625DFF7FFF86C618000003FEBE87FFFFFFFF;
defparam prom_inst_19.INIT_RAM_22 = 256'hFFFFF0C8E0100007425721FFFFFFFFFC0E60008B03FFFFFFFFFF007D10EA1F2D;
defparam prom_inst_19.INIT_RAM_23 = 256'h58006580FFFFFFFFFFE0072A83F63F02F42CFB8006240C1EAFFFEFAB58D8BFDD;
defparam prom_inst_19.INIT_RAM_24 = 256'hC3BFF201F58FA017FFFFE7F63AFEEF3FFFFC3ACC2BC007FF28303FFFFFFFFC07;
defparam prom_inst_19.INIT_RAM_25 = 256'hFF8334D55F568BA0381FFFFFFFFC00C60013602FFFFFFFFFF401C55D4446C477;
defparam prom_inst_19.INIT_RAM_26 = 256'h16D00FFFFFFFFFF80039A9F95F5FB9D877F000FE041460EFFFFFFF77FE7FFFFF;
defparam prom_inst_19.INIT_RAM_27 = 256'hF4C03B07F9C87FFFFFF7B7FFFFFFFFFFF0F5466C55737AD60FFFFFFFF88145C0;
defparam prom_inst_19.INIT_RAM_28 = 256'h0E42B9DDB737E70FFFFFFFFF0063700FCC03FFFFFFFFFFC00F146EBFB6FF8E25;
defparam prom_inst_19.INIT_RAM_29 = 256'h807FEFFFFFFC6001E65F4DF3BEFE6477C00C81FE650DFFFFFFF7FBFFBFFFFFFE;
defparam prom_inst_19.INIT_RAM_2A = 256'h8BA0FF9865AFFFFFFFFFFFFFFFFFFFC1C5CFF3F3061983FFFFFFF600200E03DB;
defparam prom_inst_19.INIT_RAM_2B = 256'h457FFEB515807FFFFDFC001D2B81C6C03FFDFFFFBFC0003CEC2E3FB745920FFC;
defparam prom_inst_19.INIT_RAM_2C = 256'h78FF7FFAE0000F8CA51F9A480EC97C01497FE33235FFFFFFFFFFFFFFFFFFF01C;
defparam prom_inst_19.INIT_RAM_2D = 256'h3FF94C0FAFFFFFFFFFFFFFFFFFFD03C6F7CAEE14C0BF7FFFE0400FCEFFF8A004;
defparam prom_inst_19.INIT_RAM_2E = 256'h8D9954C01FBFFEB8800726BDFA8C020FFDBFC6024000F9DA6CF8B0602D1780DE;
defparam prom_inst_19.INIT_RAM_2F = 256'hF9EE0300001F1DEADF9D306B9CE07B1FFCC701F7FFFFFFFFFFFFFFFFFFE03C65;
defparam prom_inst_19.INIT_RAM_30 = 256'h2109DDFFFFFFFFFFFFFFFFFFF801E39A224CE00B5CBBA81001FCAFF90300013F;
defparam prom_inst_19.INIT_RAM_31 = 256'h71E002BB9070000060B1FDFBC01019E05280000007E1958DFF27121A4835C7FE;
defparam prom_inst_19.INIT_RAM_32 = 256'hA0000000FE1B5B3F951F4A987F71FF9440330FFFFFFFFFFFFFFFFFFF401F0F00;
defparam prom_inst_19.INIT_RAM_33 = 256'h070FFFFFFFFFFFFFFFFFFFE000FC0103E0003CEC1000003C14FE7AB0000A4024;
defparam prom_inst_19.INIT_RAM_34 = 256'h000DC80400001E0D3F2F1C04122080040000000FC3352BFBB7D8BE8D0CFFCF10;
defparam prom_inst_19.INIT_RAM_35 = 256'h000000FE3B550FFB778BEF0B1FF28141187FFFFFFFFFFFFFFFFFFE000FFFFF80;
defparam prom_inst_19.INIT_RAM_36 = 256'h2FFFFFFFFFFFFFFFFFFFF0007FFF8000A40000800007029FCFE7000000000000;
defparam prom_inst_19.INIT_RAM_37 = 256'h0100200002D86FF3DDC000002000000000003FC1B76ABEC7F32326E7F180616E;
defparam prom_inst_19.INIT_RAM_38 = 256'h0003FC1AC7A0B1FD7297D87C10C0AEB1FFFFFFFFFFFFFFFFFF3E000000000408;
defparam prom_inst_19.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFECF000000000030010000000FA13FD357000000000000000;
defparam prom_inst_19.INIT_RAM_3A = 256'h0000001F79FF1C5C0000000000000000007FC1ABFA0E87A1B08E1F361012367F;
defparam prom_inst_19.INIT_RAM_3B = 256'h07FE1ADD806A34951503CD8801D35FFFFFFFFFFFFFFFF7FEBE00000002000000;
defparam prom_inst_19.INIT_RAM_3C = 256'hFFFFFFFFFFBF4E1D0000000002000000000003E3FFDEAE000000000000000000;
defparam prom_inst_19.INIT_RAM_3D = 256'h00007FFFF59BC00000000000000000007FE0A4B00EBF1BA0406381001C17FFFF;
defparam prom_inst_19.INIT_RAM_3E = 256'hFF094640FDAF44101CE20002F4FFFF7FFFFFFFFFFBF3F5800000000000000000;
defparam prom_inst_19.INIT_RAM_3F = 256'hFFFFFFF636DE780000000000000000000007F178FAC000000000000000000017;

pROM prom_inst_20 (
    .DO({prom_inst_20_dout_w[29:0],prom_inst_20_dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_20.READ_MODE = 1'b1;
defparam prom_inst_20.BIT_WIDTH = 2;
defparam prom_inst_20.RESET_MODE = "SYNC";
defparam prom_inst_20.INIT_RAM_00 = 256'hD92C4FFF3B0279F844BCCF958962F3D9621C8404D08041BEDD595A695E0671AA;
defparam prom_inst_20.INIT_RAM_01 = 256'h9550BC150CE05B51827FC100DC5095C40454000001415019055C00FAA1450EA5;
defparam prom_inst_20.INIT_RAM_02 = 256'h405451E51C7CCF083F0C1FFFEEEEBB596599B96AAA596558551F07C0D01FFE8E;
defparam prom_inst_20.INIT_RAM_03 = 256'hE0E93D1A3001B6F32C89DA69E5A05E4F6615143E62F273811555552849C95A20;
defparam prom_inst_20.INIT_RAM_04 = 256'h44001103985F38E9FCFC0455053F532174C07C7C150C500DF00FCF54530AF54B;
defparam prom_inst_20.INIT_RAM_05 = 256'h002301C01C8E8EFE010E9E4EEBB65AD99A6A5AB59C541C513FB70D323BF8FD56;
defparam prom_inst_20.INIT_RAM_06 = 256'h505C888539C7E2358FAD8200B2B6CC91F16D9A2B5E6FD7111155C45591115544;
defparam prom_inst_20.INIT_RAM_07 = 256'h06B95BC28A60FFFCC0F0D03E414E0370F4FC7C40000C00000BAAFB558BFA3E62;
defparam prom_inst_20.INIT_RAM_08 = 256'h000F03AAEAEFE7BCFEBAAAEBE6653A0449A64581000D0003A2FE0FEEEE6A1541;
defparam prom_inst_20.INIT_RAM_09 = 256'h53308D40B7F18439061A2293DAD256612C1360CB60C154499154065551455FC3;
defparam prom_inst_20.INIT_RAM_0A = 256'h54B4829C65E030FEB20303BC3EAFFFFE0037F3424C4C4CFFFAEBA980FE4B8BE4;
defparam prom_inst_20.INIT_RAM_0B = 256'h079299D78EAFEEE4AEEAA5299A6916125150D2FFCCFFEF0FCF6BEBF1A961412C;
defparam prom_inst_20.INIT_RAM_0C = 256'h3818C912FF79107E7A640A6C54190519FAC899F01571408149F0C415F004EFFC;
defparam prom_inst_20.INIT_RAM_0D = 256'hF17F06A7FEFFCFB030F383FEC3F3FFC33CCC0BF333EFFFFE8EFFA04E13897A12;
defparam prom_inst_20.INIT_RAM_0E = 256'hBD8AABBEEDA7B9AEAA51591A5154453C73EFFBDFEDEA9BAE9BFF155591265153;
defparam prom_inst_20.INIT_RAM_0F = 256'h517C41474E771E2245C0C5AD9011A510792BC030017355440D388036BDF0AEAD;
defparam prom_inst_20.INIT_RAM_10 = 256'h01569BFABEB6CDEFFECBBEBABBBFFCF3D0FB3CFFFBF3FFBF9E995792B8AAB65B;
defparam prom_inst_20.INIT_RAM_11 = 256'hA668B9ABE99D955916A1F5C9950183CFF83EEAE2A66A67EF3965543A494314FE;
defparam prom_inst_20.INIT_RAM_12 = 256'hDAB843CC5ECC7DCBEA8A2E83D5AFE696EC033C17149645331CBC702AEABEC670;
defparam prom_inst_20.INIT_RAM_13 = 256'h55E5E956ABB6ABCF6AA9AEDAFEBFBC33F0EBAFFB4FF3F3AF9A13A4B97E307F35;
defparam prom_inst_20.INIT_RAM_14 = 256'hB56D557899811451C6154043CE2CBBBEBA3B85A695AAE995994496011040D519;
defparam prom_inst_20.INIT_RAM_15 = 256'h52B11201B4C776A85564CB7FC15EDBFCFCC134084C33CF3CF33AA5B964230542;
defparam prom_inst_20.INIT_RAM_16 = 256'hAAAAAAAA659EAF59A795BBAA6AAF70F3FEAAFBFF3000FBEE53919836487ED0E9;
defparam prom_inst_20.INIT_RAM_17 = 256'hA5952A9450D355810410AFFAD6FAAA525559645696A4C5445584110443556554;
defparam prom_inst_20.INIT_RAM_18 = 256'h4CCCA3ABE924965E5DA280FD41EEFC0342CF3C3FF32F3F4AA2B5A99972695959;
defparam prom_inst_20.INIT_RAM_19 = 256'hE152E0650A859AA156BAFA6E96BBEEFBEAF2060F0CFF5A82D49B02CCC4D49831;
defparam prom_inst_20.INIT_RAM_1A = 256'h444043140943C00CC7BFAA9979413E51112956A21455017DC5105551515A551A;
defparam prom_inst_20.INIT_RAM_1B = 256'h651EF91ABD68108B08EE5F46FFCFAFFCF3FFEA6471B3A8E8A665059140552744;
defparam prom_inst_20.INIT_RAM_1C = 256'h45C55216505415525259AAA76E76BAA0E0C04010FE8653E35782B5701D44D9A7;
defparam prom_inst_20.INIT_RAM_1D = 256'hC42C3C7483C030FBA400740F31E471110444854550147479000585855D46A475;
defparam prom_inst_20.INIT_RAM_1E = 256'hF6360FB9821E441CAEF1A5FEEAFEC26F3ABED1AA96669591B400C400CC544501;
defparam prom_inst_20.INIT_RAM_1F = 256'h5551654183F5411574AABAA969EBAB3CF041CC3FF3909232AF675C86C2BDDC72;
defparam prom_inst_20.INIT_RAM_20 = 256'h03690CFFDF62E157442F0033043F071F500C100002FF0001545409F4535516C0;
defparam prom_inst_20.INIT_RAM_21 = 256'h470C7363F1FF611AD4A9F77F6AABA28B1B179A6A5455800333FCEF13007C0F3C;
defparam prom_inst_20.INIT_RAM_22 = 256'h31730E014180D55448952A9AF3E00F00547443BA8F5E2FFBF9924138C9629D21;
defparam prom_inst_20.INIT_RAM_23 = 256'h64FBCE8EF95D0573FB2394CA08CDD31CC3D3CFFEBCC0F213FFC0F35FF31F10D3;
defparam prom_inst_20.INIT_RAM_24 = 256'h7922C8F1186586AAAABA96982FE9AAAF95A290F6B6CCBEEEB1D3C3EFE8F0C0E3;
defparam prom_inst_20.INIT_RAM_25 = 256'h0B3F3C0003D405595959A8EC000005374440FF9389F7E16313C1529658A0B1F7;
defparam prom_inst_20.INIT_RAM_26 = 256'hF3BEEE5040FFF0BFEE8FFA3BBDBCBBFF3FBFD3C104C4F0F00FCF5F0CF00C733F;
defparam prom_inst_20.INIT_RAM_27 = 256'h3B72D6A29F2516A9A95B6AB9ED571428663CFF0333F6EFFABC23828BBBEFEFBB;
defparam prom_inst_20.INIT_RAM_28 = 256'hEFF0FEB8350445555AAAAA3015A1095003355F8B811FF8C63CF5F419E3011DED;
defparam prom_inst_20.INIT_RAM_29 = 256'hE66D3804BBAEFD93A9FFCF0FBF3B23BF2EE2F0EE3BEBB0FFCFFCFF2FEC4EBF4E;
defparam prom_inst_20.INIT_RAM_2A = 256'h741452F08165E51DA1EB9AE1B5D0603E7FDC1ABA29B5BFEFEBFBF3FBD73ABBBF;
defparam prom_inst_20.INIT_RAM_2B = 256'hD63FBE01015955A80AA400552A950287E972B0635065549FA4AF9F04310773D9;
defparam prom_inst_20.INIT_RAM_2C = 256'hCBBEF619DFDF66A6995AABFAFBB947FBEFFF6BBEC08FFDA2BF0CAF9ADFEA27AA;
defparam prom_inst_20.INIT_RAM_2D = 256'h609F025A6AA97229954A961428C8E4D7FBFD771A5ABAD2B59761EE332AB6A5A4;
defparam prom_inst_20.INIT_RAM_2E = 256'h9723FCF0C01956AB8C00025055824CF90E23339EF8DCC9489781ECCEB5257635;
defparam prom_inst_20.INIT_RAM_2F = 256'hF6AE1580496AE449A9856BEAAA6C587BA3BBBEFAAFF2A4BABA8F8A9AAAAAABEE;
defparam prom_inst_20.INIT_RAM_30 = 256'h81111554541044E50457FE60B6EA62AA456F945A5299B26ACADA25A94AA4A70F;
defparam prom_inst_20.INIT_RAM_31 = 256'hBFF0CFF05657038C50175AA6A803E60E22153FCDD5D681ED07BD038D50ADA3C6;
defparam prom_inst_20.INIT_RAM_32 = 256'hA565A5654636A43B5525AA9684292B2D7A6AAE5B1B428E2AA86956A12A956BE7;
defparam prom_inst_20.INIT_RAM_33 = 256'h543550113100940B76EA9F752759567556924866745084656355A12C033BA956;
defparam prom_inst_20.INIT_RAM_34 = 256'h7BF555C56A4BC041D5456A9542EA75A106201A97B73843DE894ED5E6F7F87C29;
defparam prom_inst_20.INIT_RAM_35 = 256'h5C56144003681965595559251568848B1560624A26525566559611555556CBEA;
defparam prom_inst_20.INIT_RAM_36 = 256'h14810010D059467397A8559505A20142225D1144005115C6600D40E666258A51;
defparam prom_inst_20.INIT_RAM_37 = 256'hC60C45F6BF3055E9596AA560A40AE2DCA4FC3F79E0D35C4479AB90F616FD9400;
defparam prom_inst_20.INIT_RAM_38 = 256'hD7C37C00C01555066DA045276851864114C0157955D401500543951546929BF2;
defparam prom_inst_20.INIT_RAM_39 = 256'h0014C161E0F75CC9425010503403981135101468300037408CED5D457F052561;
defparam prom_inst_20.INIT_RAM_3A = 256'h5146ABB0105A2AA295A5D3AAC4ED2BC6E9A01CF938AFAB1F878073AC134013B2;
defparam prom_inst_20.INIT_RAM_3B = 256'hC0CF4F72F873CC8C10D4989111D074B73EC00511D0103050FDB0144955857B40;
defparam prom_inst_20.INIT_RAM_3C = 256'h240E0DC8CA9D4FF1B159101436678C01D241CDF008ED0FBBC54451EB832F4EED;
defparam prom_inst_20.INIT_RAM_3D = 256'h0AEB0C0045A9ABDA550FF2E5D9BD6B16E1D9A16A075CB02CCB052D1410DFB3D0;
defparam prom_inst_20.INIT_RAM_3E = 256'hF653303CE30D410C0009C0C400333CF5F133053FFCEFC3CF000500165ABBBFC1;
defparam prom_inst_20.INIT_RAM_3F = 256'h7CEC61F08C2AD0FC5F1F9F103FFFBFBFFFB7FB8FFFA6929705102CC003EAFC3C;

pROM prom_inst_21 (
    .DO({prom_inst_21_dout_w[29:0],prom_inst_21_dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_21.READ_MODE = 1'b1;
defparam prom_inst_21.BIT_WIDTH = 2;
defparam prom_inst_21.RESET_MODE = "SYNC";
defparam prom_inst_21.INIT_RAM_00 = 256'hAA90E3B16D5540EE5D4CCC60D5AC596A49D151551500FAA916AAAAAAA6AAAAAA;
defparam prom_inst_21.INIT_RAM_01 = 256'h0000FC000CFE2FCA7F0015551155551555555555555555555551550000000FFF;
defparam prom_inst_21.INIT_RAM_02 = 256'hAAAAAA9AA69665A695A6A5555555555555555555555555555550541515500010;
defparam prom_inst_21.INIT_RAM_03 = 256'h54E4C1ED7554EECB0C15E21BB15A93DC6255554002AB256AAAAAAAAAAABAAAAA;
defparam prom_inst_21.INIT_RAM_04 = 256'h00000003E4ABCBC00101555555405455451541415551555105501000030FFFFA;
defparam prom_inst_21.INIT_RAM_05 = 256'hAAA9AA6A96656555AAA555655555555555555555515551554004514440010000;
defparam prom_inst_21.INIT_RAM_06 = 256'h39C26E9140FEE330D4786EC5992712C45541003E7F1569AAAAAAAAAAAAAAAAAA;
defparam prom_inst_21.INIT_RAM_07 = 256'h00300FA146F0000115051541555154450501415555515555500000000FFFEA94;
defparam prom_inst_21.INIT_RAM_08 = 256'hAAA5A95555555956555555555555555555555555555155540400500000000000;
defparam prom_inst_21.INIT_RAM_09 = 256'hC1AED154F17B0F3DF2AA1950305555554143E7C15A6AAAAAAAAAAAAAAAAAA569;
defparam prom_inst_21.INIT_RAM_0A = 256'h00FFAABC000545000454540140000000554404545151510000000000FFFAA4F9;
defparam prom_inst_21.INIT_RAM_0B = 256'hA55965556555555555555555555555555555150011000050100000000000000C;
defparam prom_inst_21.INIT_RAM_0C = 256'h9A95103E92E3DCFDAC54A32655555500FF8C155AAA9AAAAAAA5A6AAA5AAA5556;
defparam prom_inst_21.INIT_RAM_0D = 256'hFFFF000000001005450414001404001441115004440000001000000FFEA538F1;
defparam prom_inst_21.INIT_RAM_0E = 256'h5555555555555555555555555555554144000000000000001000400000000003;
defparam prom_inst_21.INIT_RAM_0F = 256'hD540F94F33FB1FF03D3C1551554403E031556A9AAA9AAAAAA6966A99565A5555;
defparam prom_inst_21.INIT_RAM_10 = 256'h000000300000100000100000000001041500410000040000000003FE9538AD99;
defparam prom_inst_21.INIT_RAM_11 = 256'h55565555555555555555151555551410014000000000000040000030000300FF;
defparam prom_inst_21.INIT_RAM_12 = 256'h00C63C59ACBAAD136155515400F8C81556A996A9AAAAAA99A6569A9555555555;
defparam prom_inst_21.INIT_RAM_13 = 256'h0000000000000010000000000000014405000000500404000003FF9534AD8A05;
defparam prom_inst_21.INIT_RAM_14 = 256'h555555455555555515555554104100000000000000000000000000000000C000;
defparam prom_inst_21.INIT_RAM_15 = 256'h77D532C1791782155555102FF7C01556566A9AA6A69965965995555556545555;
defparam prom_inst_21.INIT_RAM_16 = 256'h00000000000000000000000000000504000000004555000003FEA528A98B1503;
defparam prom_inst_21.INIT_RAM_17 = 256'h55555555555455555555000000000000000000000000C0000000000003000000;
defparam prom_inst_21.INIT_RAM_18 = 256'h404AC4039D3155515004F80C155556A9A9659695599595555955555545555555;
defparam prom_inst_21.INIT_RAM_19 = 256'h000000000000000000000000000000000004545051000003FFA437699D150E85;
defparam prom_inst_21.INIT_RAM_1A = 256'h55555555555415511400000000003C00000000000000003CC000000000000000;
defparam prom_inst_21.INIT_RAM_1B = 256'hAC0D4600B15515031B1EC0555565555659555556595955555555555555555555;
defparam prom_inst_21.INIT_RAM_1C = 256'h00C0000000000000000000000000000505155555001003FEA4F709BF50085203;
defparam prom_inst_21.INIT_RAM_1D = 256'h15514145141545000000300F30C030000000000000003030000000000C000030;
defparam prom_inst_21.INIT_RAM_1E = 256'h154051C55540067D7C0555555555699595555555555555554555155511555555;
defparam prom_inst_21.INIT_RAM_1F = 256'h00000000C3F000003000000000000041055511400400FE94E2048D14210E70AA;
defparam prom_inst_21.INIT_RAM_20 = 256'h5441510010440003000F0033003F030F000C000003FF0000000000F0030000C0;
defparam prom_inst_21.INIT_RAM_21 = 256'h5450444703F9B700155555955555596595955555555555544401005455415041;
defparam prom_inst_21.INIT_RAM_22 = 256'h30330F000000C0000000000004055055554554000FFA9392C58D53FA70F77A45;
defparam prom_inst_21.INIT_RAM_23 = 256'h05001010000C0033FF33C0CC0CCCC30CC3C3CFFFFCC0F003FFC0F30FF30F00C3;
defparam prom_inst_21.INIT_RAM_24 = 256'h3D4410338DB01555555555565555555455555504051100000404140001051504;
defparam prom_inst_21.INIT_RAM_25 = 256'h0F3F3C0003C00000000001015555554455550003FA4392C9AC54FD7F0CAA4504;
defparam prom_inst_21.INIT_RAM_26 = 256'h0400000000FFF0FFFFCFFF3FFCFCFFFF3FFFC3C000C0F0F00FCF0F0CF00C333F;
defparam prom_inst_21.INIT_RAM_27 = 256'h0033FA8F00555555555555555555555655410054440000000144141000000000;
defparam prom_inst_21.INIT_RAM_28 = 256'hFFF0FFFC30000000000000455555555554400FF9539DCA6E3B67E83A545551C0;
defparam prom_inst_21.INIT_RAM_29 = 256'h000C3C0CFFFFFFF3FFFFCF0FFF3F33FF3FF3F0FF3FFFF0FFCFFCFF3FFC0FFF0F;
defparam prom_inst_21.INIT_RAM_2A = 256'h3E2EC00555555555555555554555554000114000400000000000040000400000;
defparam prom_inst_21.INIT_RAM_2B = 256'hCF3FFF000000000000015555555555540033EA428EDC8297C6EFA55545433000;
defparam prom_inst_21.INIT_RAM_2C = 256'hCFFFFF3CFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFC0CFFFF3FF0CFFFFCFFF3FFF;
defparam prom_inst_21.INIT_RAM_2D = 256'hAC00555555555555555555554111010000000000003000000000000440300000;
defparam prom_inst_21.INIT_RAM_2E = 256'hFF33FCF0C000000011555555555551000FE94249DD4B8B96E9551110040033C2;
defparam prom_inst_21.INIT_RAM_2F = 256'hFFFFFFF3FFFFFFFFFFCFFFFFFFFCFCFFF3FFFFFFFFFFFCFFFFCFCFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_30 = 256'h155555555555555555540005000004000000000000000000000000000000330F;
defparam prom_inst_21.INIT_RAM_31 = 256'hFFF0CFF000005411555455555554000FE94E78EC560166F15400018000EBBAC0;
defparam prom_inst_21.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF3FFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_33 = 256'h5545555545555554440000300000003000000000000000000000000C033FFFFF;
defparam prom_inst_21.INIT_RAM_34 = 256'hFFF000C0001015551555555554003FA94E7933399E9B3010029730FCD5BC0155;
defparam prom_inst_21.INIT_RAM_35 = 256'hFFFFFFFFFEFFFFFFFFFFFBFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_36 = 256'h55555555155154440300000000030000000C0000000000C0000C00FFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_37 = 256'hC30C00000045551555555555000FA93A7A2E973FBD30355CFEFE036F00015555;
defparam prom_inst_21.INIT_RAM_38 = 256'hBEBEEBFFBFFFFFFFFBFFFFFEFFFFFFFFFFBFFFFFFFBFFFFFFFFEFFFFFFFFFFF3;
defparam prom_inst_21.INIT_RAM_39 = 256'h554515450504000003000000300300003000003030003300CCFFFFFFEAFFFFFF;
defparam prom_inst_21.INIT_RAM_3A = 256'h000000055551555555551400CFA5390E29F9E8D6AFBBEABA90BBF00154555445;
defparam prom_inst_21.INIT_RAM_3B = 256'hBFBAFAEEABEEBBFBFFBFFFFFFFBFEFEEEBBFFFFFBFFFEFFFABAFFFFFFFFFFFC0;
defparam prom_inst_21.INIT_RAM_3C = 256'h45505111100C0FF0300C30003333CC00C300CCF00CCC0FFFFFFFFFAEFEEAFAAA;
defparam prom_inst_21.INIT_RAM_3D = 256'h0000515555555555555000FFA53A4D1B374390FDB9640372BF01415555100415;
defparam prom_inst_21.INIT_RAM_3E = 256'hAEBEEFEBBEFBFFFBFFFFBFBFFFEEEBAFAFEEFFEAABAABEBAFFFFFFFFFFFFFFC0;
defparam prom_inst_21.INIT_RAM_3F = 256'h41010500CC3FC0FCCE3FFF303FFFFFFFFFFFFFCFFFFFFFFEFFFFEBBFFEAAABEB;

pROM prom_inst_22 (
    .DO({prom_inst_22_dout_w[27:0],prom_inst_22_dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_8),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_22.READ_MODE = 1'b1;
defparam prom_inst_22.BIT_WIDTH = 4;
defparam prom_inst_22.RESET_MODE = "SYNC";
defparam prom_inst_22.INIT_RAM_00 = 256'hFDE33D3937578774455AD22E68CCF00214344345432444434444335133431335;
defparam prom_inst_22.INIT_RAM_01 = 256'h11223433345655666677666666555564443323220ECB98642FB992D5E702C751;
defparam prom_inst_22.INIT_RAM_02 = 256'hBBBBCCBBBABABBCBCB9ACBCBABBCCBBCBBCBBDBCBCCEDCCEEEDFEFF000112232;
defparam prom_inst_22.INIT_RAM_03 = 256'hBAA9CBBBBBBCCBBBCBBBBCCCBACCCBBDBACCACBBCABBABCBCBBBBBCCADBBBACB;
defparam prom_inst_22.INIT_RAM_04 = 256'hEECEEF0EF0FE0EFEECBCCCDDCBCBBCABCAAAA9AB9AACB9B9AACACBBAABBBBCAB;
defparam prom_inst_22.INIT_RAM_05 = 256'h5233103302011F0FEEF00FFEEFEEEEFFEDDEFFEEFEEEEEFFFEEFEEEFFFEF0EEE;
defparam prom_inst_22.INIT_RAM_06 = 256'h0B08CA84FF2E4645C39AC0003244423533525443334336134144324444233131;
defparam prom_inst_22.INIT_RAM_07 = 256'h4253454436675766657566665545443322010EFCB9952FB972C51A143D9F659E;
defparam prom_inst_22.INIT_RAM_08 = 256'hBBBA99ACABBB9AC9ABCCABBAABAABCACCBCCCDDDCEFFFCFEF00002F123214234;
defparam prom_inst_22.INIT_RAM_09 = 256'hAABCDBBAAADCCABCABBABBCBCB8CBCDBAA9AABABCCCBBBBBCCADAA99BBBABCAA;
defparam prom_inst_22.INIT_RAM_0A = 256'hD0DDEEEDFCDCECBCBBCBBBCAA9ABBA89ABABAA8BBABA8ABAAAABA99BEAA889AA;
defparam prom_inst_22.INIT_RAM_0B = 256'h110F00FEEFEDEEEFCE1EDFFFFFFFFFECEDEFDDDEFCCDFDDDCCCCFEDEDDDFDDD0;
defparam prom_inst_22.INIT_RAM_0C = 256'h075EE8983B88ACDFF02333444454443434333242242333134413323221241131;
defparam prom_inst_22.INIT_RAM_0D = 256'h5554565663666665565665554442200FEEEBA87542F961D71A3F9E776BE032FF;
defparam prom_inst_22.INIT_RAM_0E = 256'h8AAA99AAA9AAAAAA9AABBBDBBBBAACBCCCDDCDDDEEEFFF001211112222234333;
defparam prom_inst_22.INIT_RAM_0F = 256'hAABAACBAABBABBBBBAACAAAA99BBBAAAAAAAAA9AA9ABAABB8A99B9A9ABAABAA9;
defparam prom_inst_22.INIT_RAM_10 = 256'hCDCBEDCBBCBBBCAAB99BB9ABAA9899999AAA99999A89ABAA9CAB9998BAAAAA8B;
defparam prom_inst_22.INIT_RAM_11 = 256'hFEFBCCECFDEEDFF10DFFCDDEEDDEEDEDEDEDDDCCCCBDEDEDDDECDDDEEBEEEDED;
defparam prom_inst_22.INIT_RAM_12 = 256'h42F588CFF0012034344544544414443322332222213112122132302120F1FF0F;
defparam prom_inst_22.INIT_RAM_13 = 256'h54668767766566666654533223011EDCC997420E750B83E857D21111234566CD;
defparam prom_inst_22.INIT_RAM_14 = 256'h7999AAAAAAA9ABBAAABABBBAAC9BCCCDDDEEEFE0FFFF01122222222323445556;
defparam prom_inst_22.INIT_RAM_15 = 256'h9CB99AAAA9AAAB9BBAB99AA7AAA99AAA99AAA9A9AB7AA998AAB8AA98AA99ABA9;
defparam prom_inst_22.INIT_RAM_16 = 256'hCCB9ABBBAAA97AA999AA9A9AAB9A99987998899BAAAAA9BAA999A9A9A98AC9A9;
defparam prom_inst_22.INIT_RAM_17 = 256'hCDEDDDDEDDEFDDDEDEDEFCDBDCCCDEDDDDCCCCDCBDDCEEBDDBCDCCECDECBCEAB;
defparam prom_inst_22.INIT_RAM_18 = 256'hEF0F0213343244442442523433342231122313322111211110200F1DE0DEEDCC;
defparam prom_inst_22.INIT_RAM_19 = 256'h67766666666654544442222010DEBB78862FBB760EC63DDDF073792319E375AB;
defparam prom_inst_22.INIT_RAM_1A = 256'h89999989AAA999AAAABAABBBBCCBCEDEDEEEE0010F2211222342345553467667;
defparam prom_inst_22.INIT_RAM_1B = 256'hA979999AA9999A9AA9999A9AA8998898898798A99B89A9998987889A98877899;
defparam prom_inst_22.INIT_RAM_1C = 256'hB9A8989989A8A89898998999789888899A988898A9989889A9A999A9A999BAA9;
defparam prom_inst_22.INIT_RAM_1D = 256'hCEDDDECCCDCDCDCDCEDBDDDCCDDDABBCCCBCBCBDADDEFCBCDBCDDDBABAA989AB;
defparam prom_inst_22.INIT_RAM_1E = 256'h3332344442252333333343322022332101F1222122101010DFEEEDDDCCCDCDCC;
defparam prom_inst_22.INIT_RAM_1F = 256'h6677566565456353422110FECCA8775430FDA8523101678CDF23568CCEE00213;
defparam prom_inst_22.INIT_RAM_20 = 256'h889A88898A999AAAACACBCCDCCDDDDE0F0F00110012424334346354565576666;
defparam prom_inst_22.INIT_RAM_21 = 256'h979988A98898997999AA8788888A88979789998798899878A677777987888988;
defparam prom_inst_22.INIT_RAM_22 = 256'h9979767897887977888897677875876778789889899899988899789899AAA9A7;
defparam prom_inst_22.INIT_RAM_23 = 256'hEDDCBCCEBDDBCBCBCACACDCCABCDABBCCABAAADBBCBABA8BAABA988989989878;
defparam prom_inst_22.INIT_RAM_24 = 256'h332333432332222131121241211110111112F0011EEEECEEFDDACCBBEECDCADD;
defparam prom_inst_22.INIT_RAM_25 = 256'h7665555455534320F0F0DECB8877432221EDECEF2305678BDEFFF11221233545;
defparam prom_inst_22.INIT_RAM_26 = 256'h79789988BBBBAABCBCCCBEFDEEFFF00000132113233362543554456666566545;
defparam prom_inst_22.INIT_RAM_27 = 256'h788798888779779898698A967887769777885887876767766578768877689888;
defparam prom_inst_22.INIT_RAM_28 = 256'h756986676787898867887887777776878778887799978B588989A77898887988;
defparam prom_inst_22.INIT_RAM_29 = 256'hBCCDBCCCDACBCCABABBA9ABD9CB9CBCCBCD9AAAAB98978897778878786888679;
defparam prom_inst_22.INIT_RAM_2A = 256'h223332222111112F1121110000012F21FEDEECECDFCCBBCB9BAABABDA9BBCBDA;
defparam prom_inst_22.INIT_RAM_2B = 256'h5455534444313110FDDCBAA887766555557679899ADE00F13222344433432222;
defparam prom_inst_22.INIT_RAM_2C = 256'h88AA9999AB9ABBADDDEEEFEFEE00000202222333343555565665666556666665;
defparam prom_inst_22.INIT_RAM_2D = 256'h7887577898779689887887775686757886665556655566767768778668878788;
defparam prom_inst_22.INIT_RAM_2E = 256'h5676776778666466766686687567877688788878779867787878885988877777;
defparam prom_inst_22.INIT_RAM_2F = 256'hA9CAACBAA9A989A7AA9A9B9AB9AAB99B88A87877777766856766745565686866;
defparam prom_inst_22.INIT_RAM_30 = 256'h2122212212112010000110F0FEDEEECDBCDDBCBBCB9B9AACBBBEBBBABBBBBCAA;
defparam prom_inst_22.INIT_RAM_31 = 256'h444433323110EFDDECBBABA9BCA9ABBADDEEFFFF312334333332323312222003;
defparam prom_inst_22.INIT_RAM_32 = 256'h89A989BBAABCCDDEDDE0000F0011222222333444454555554655665665555445;
defparam prom_inst_22.INIT_RAM_33 = 256'h7867776674656556667667656665456554545655567557665676675776669989;
defparam prom_inst_22.INIT_RAM_34 = 256'h5565757655667668867665675776766688665876667667676686676787886777;
defparam prom_inst_22.INIT_RAM_35 = 256'h9B9999A98999989AAA8A99AA9A87777655576455655666656654565656437566;
defparam prom_inst_22.INIT_RAM_36 = 256'h00000000000000000000000000000000A9BB999BA8AA9AAAAA99BBABBB98A898;

pROM prom_inst_23 (
    .DO({prom_inst_23_dout_w[30:0],prom_inst_23_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_23.READ_MODE = 1'b1;
defparam prom_inst_23.BIT_WIDTH = 1;
defparam prom_inst_23.RESET_MODE = "SYNC";
defparam prom_inst_23.INIT_RAM_00 = 256'h0000000931EDFFFFFFFFFFFFFFFFBFFFFFFF679FFFFFFFFFFFFFFFFFFFFFFFFA;
defparam prom_inst_23.INIT_RAM_01 = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFB800000;
defparam prom_inst_23.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFF600000000000000403F7EFFFF767FFDFF87DBFFFF;
defparam prom_inst_23.INIT_RAM_03 = 256'h000021597FFFFFFFFFFFFCFFBA7FFFFFDC6DBFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_04 = 256'hE7DDD7FFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFE1000005000;
defparam prom_inst_23.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFEC000006F8000000001397DFFF9FFFFFFC819F61D8007;
defparam prom_inst_23.INIT_RAM_06 = 256'h0000184EF7FE79FFFF300210006001999A76FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_07 = 256'hE0FCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFED000002FF80000;
defparam prom_inst_23.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFBE4000002FFFE0000000021B79DFFFFF4C0208100108032B43;
defparam prom_inst_23.INIT_RAM_09 = 256'h0100637FB41E8600000040400B664A2D02CFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0A = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB208000057FFF4000000;
defparam prom_inst_23.INIT_RAM_0B = 256'hFFFFFFFFFFEF42000017FFFEC00000005818FFE807A0800008205002C86A8860;
defparam prom_inst_23.INIT_RAM_0C = 256'h01FF8696003008200000001049C0027FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7400000DFFFF6F00000000;
defparam prom_inst_23.INIT_RAM_0E = 256'hFFFFFFFFFB0000079FFF77A0000108007FE020800C0100000000001A800037FF;
defparam prom_inst_23.INIT_RAM_0F = 256'hFE068000000200000000184E081FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF340000A39FF39F6000000241F;
defparam prom_inst_23.INIT_RAM_11 = 256'hFFFFFD008003E3CFB9FF3000100539F786440C000000002000038AEF0DFCFFFF;
defparam prom_inst_23.INIT_RAM_12 = 256'h910300000000000000622DC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBB40400FFE39D8FFF2A04100CFFBE1;
defparam prom_inst_23.INIT_RAM_14 = 256'hFFA4000FFFEBFDFFFFA007F9FE7FDB837000000000001080009D1C73FFFFFFFF;
defparam prom_inst_23.INIT_RAM_15 = 256'h10000C000008000001844F5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000EFFFE30FFFFED3FF7DFFFFDF962;
defparam prom_inst_23.INIT_RAM_17 = 256'h8002FFFFFDDFFFE6BFFFFFFFFEEFF88000F000000000000042EC5FEFFFEFEFFF;
defparam prom_inst_23.INIT_RAM_18 = 256'h0240018100000000F8FFFDFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_23.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB68057FFFCF9DFFFF3FFFFFFFEFFF7A0000;
defparam prom_inst_23.INIT_RAM_1A = 256'hEFFFEE71DFF33FFFFFEFFFFFE6C00000000068400000602233FFFFBFFFBFFFFF;
defparam prom_inst_23.INIT_RAM_1B = 256'h0000800000003D3FDAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC400;
defparam prom_inst_23.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFBF1272E7FEF3F1FFB9FFFFDFFFFFFFE60000000;
defparam prom_inst_23.INIT_RAM_1D = 256'hFF3FE1F99FFFFBFFFFFFFFE00000000101010000000B0EFFCFFFFFFF7FFFFFFF;
defparam prom_inst_23.INIT_RAM_1E = 256'hC0A0000002C3FFDFDFEFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEB603C67;
defparam prom_inst_23.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFBF1FF8E73BFFF5FDFFFFFFFFFFFFFF8000000FF01;
defparam prom_inst_23.INIT_RAM_20 = 256'hFFFDC7FFFEDFFFFFFF7618000BFA91400055002020FFAFFFF7FFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_21 = 256'h0100004F97DFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFCBFF8EF8F;
defparam prom_inst_23.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFBFDFFF87CFFFFC96FFFE6FFFFFFFF4800005F3DF8200;
defparam prom_inst_23.INIT_RAM_23 = 256'h69EFFF6FFFFFFFF6400001EF77BC000025010307FBFFFBFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_24 = 256'h40016FDFDBFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBDFFFFE7FFFFC;
defparam prom_inst_23.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFF3EFFFFCD7FFFEF7DFFF737FFFFFFF400003DC06BD800000;
defparam prom_inst_23.INIT_RAM_26 = 256'hFFBFDFFFFFFE480003CFAA06E00000100269F7F9FBFDFFEFFFF7FFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_27 = 256'h000FFDFFF77B3FE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCDBFFFCE7FFFE33FD;
defparam prom_inst_23.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFEB3FFE662FFE38FF5F18FFFFFFFFF000206B13CA7E00000400;
defparam prom_inst_23.INIT_RAM_29 = 256'hFFFFFFFFFC80003BA80E0C60000000000EDFFFBCFCD97FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2A = 256'h87FFFF3F33DFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB3FEE5FE799CFFF0FC;
defparam prom_inst_23.INIT_RAM_2B = 256'hFFFFFFFFFFFF43BEF1FFE79CFFFF0F7FFFFFFFFD20001FFBC62FFE0000000003;
defparam prom_inst_23.INIT_RAM_2C = 256'hFFFFFFA000079F28BFFF90000000001EEFFE7FF7B9FFFBFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2D = 256'hF3FFFFBFEEDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEB379FFFE7E7FFFE0BFDF;
defparam prom_inst_23.INIT_RAM_2E = 256'hFFFFFFFFFDEBB8FFFF668FFFF3BFF7FFFFFFD60043F3F0FFFFBC00000000003C;
defparam prom_inst_23.INIT_RAM_2F = 256'hFFE60200FE7CFFFFEF00000000000C3E7FDBDDFBF1FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_30 = 256'hB7FEFFEEFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBCFFFF87BBFFFF57FFFFFF;
defparam prom_inst_23.INIT_RAM_31 = 256'hFFFFFFEFF4FFFFCF273FFBB4FFFFFFFFFD40003FCF7FFF33F00000000000BF3F;
defparam prom_inst_23.INIT_RAM_32 = 256'hD0203FF9DFFEE57D00005880001FCFFFE6BEFBDFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_33 = 256'h9EFE7FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFBFDF7FFF30E7BFDAF3F7FFFFFFF;
defparam prom_inst_23.INIT_RAM_34 = 256'hFFFF7FC7FFD78E673CCFDF9FFFFFFFF800017F1FFDD82F80001DEA01004DFFFB;
defparam prom_inst_23.INIT_RAM_35 = 256'h0017C7FF0C03F80008001080C3EEF597FCFFFEFFFBFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_36 = 256'h6167FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE67FF3CFF6767FE7CBFFFFFFFFC0;
defparam prom_inst_23.INIT_RAM_37 = 256'hF7FEE7FBC7FE67E7F9EF3FFFFFFFF00047FAFF09483E000580062433F8BFE3FE;
defparam prom_inst_23.INIT_RAM_38 = 256'hFF7C004027A00026020026DCFDFBF7FCDF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_39 = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFE7E9CF9E7FFFB73FE05EFFFFFFDDC284F;
defparam prom_inst_23.INIT_RAM_3A = 256'hC7CFE3DFFE29FFC3F3FFFFFFFF5D73FFCF200341F80000002001A37FFF4FFFAF;
defparam prom_inst_23.INIT_RAM_3B = 256'h9C60402F000000002037FFEFE77FA7E76B3FFFFFFFFFFFFFFFFFFFFFFFFFFFE7;
defparam prom_inst_23.INIT_RAM_3C = 256'hFDFFFFFFFFFFFFFFFFFFFFFFFFFFF77FFEF3FFBFBB7FF27E7FFFFFFFFFDDFFF9;
defparam prom_inst_23.INIT_RAM_3D = 256'hC30FFFCBBFFD7F04FFFFFFFFFFFFFF94810C41F00000000058CCFFFE19E76E1B;
defparam prom_inst_23.INIT_RAM_3E = 256'h01007C0000000026333FFF9E79D9E3FF7FFFFFFFFFFFFFFFFFFFFFFFFFFC773F;
defparam prom_inst_23.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7F1FFD77FFCDC7FDDFF0FFFFFFFFFFFFFFF110;

pROM prom_inst_24 (
    .DO({prom_inst_24_dout_w[30:0],prom_inst_24_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_24.READ_MODE = 1'b1;
defparam prom_inst_24.BIT_WIDTH = 1;
defparam prom_inst_24.RESET_MODE = "SYNC";
defparam prom_inst_24.INIT_RAM_00 = 256'hBFE572FDCFF40FFFFFFFFFF2FFFF2E02115FC00000800B40FEF5F87E4423314F;
defparam prom_inst_24.INIT_RAM_01 = 256'h02F00000000037FEFFBFE7E3F93D77FFFFFFFFFFFFFFFFFFFFFFFFFFEBF3FEF7;
defparam prom_inst_24.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE7FFBD73CE3EFE57FC01FFFFFFFF9B7DFFF1C20E;
defparam prom_inst_24.INIT_RAM_03 = 256'h3FEE2CFF007FFFFFFFEFADDFFEF800097F0000000004FF9FEB79F167BEFF6FFF;
defparam prom_inst_24.INIT_RAM_04 = 256'hE0000000848EBDFFFFF03877DFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEFFDD737;
defparam prom_inst_24.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFE4FDFD7F5FFFBF3F201FFFFFFF5D26A83FCE041C07;
defparam prom_inst_24.INIT_RAM_06 = 256'hD3CF0007FFFFFE9B4F33F7F98008137E00000002236F779F7B873FF9FFFFFFFF;
defparam prom_inst_24.INIT_RAM_07 = 256'h000000015FFFDEFE40817EFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F8FD7FD7BFF4;
defparam prom_inst_24.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFF33FBFD1FFF4BE3F503FFFFFEFAFBDF265F2010246FE0;
defparam prom_inst_24.INIT_RAM_09 = 256'hC441FFFFFEF7E09DEDA5E4086C0BFC000000003FFDFFFFF967FFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0A = 256'h000C3FFFFFFFE6187FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDF86B9FFEFFF0BF8;
defparam prom_inst_24.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFDFBE3DFFFFFC7FE32107FFFFF7ED901FF94FC8018105F8000;
defparam prom_inst_24.INIT_RAM_0C = 256'h3FFFFF9ED5C0CD76EF9020300BF02000002DFFFFF8E011F978DEFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0D = 256'h13FFDF9E7F1AED1FFF7FFFFFFFFFFFFFFFFFFFF7FFFFFD9E7F3FFDFFE17F8264;
defparam prom_inst_24.INIT_RAM_0E = 256'hFFFF7FFFFFFFF94FE2FFFFFA5FE1B11FFFFFCFA90C036DCFF204A1107F400100;
defparam prom_inst_24.INIT_RAM_0F = 256'hFFE5D91FFE1A363E48C8C01FF00000009FF7FFDF9F78A7EFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_10 = 256'hDFFFFDE7A0F8DDFFFFFFFFFFFFFFFFEFFF9FFFB7FFDFA3FCBFFFF1D7E0DC47FF;
defparam prom_inst_24.INIT_RAM_11 = 256'hEFEFBF7FF7F8FFA1F97A2FFD9F0FFFFFF1899FFFF0B757CB010091FFFB0003DF;
defparam prom_inst_24.INIT_RAM_12 = 256'h63CFFFFF89F9796381807FFE4200FFF4FFFEFFF90F375FFFFFFFFFFFFFFFFBFF;
defparam prom_inst_24.INIT_RAM_13 = 256'hFFFFF3847F7DFFFFFFFFFFFFFFFFFEFF1BFFDFFDFD9FFC3F5C7B7C6799FFFFFC;
defparam prom_inst_24.INIT_RAM_14 = 256'hFB3FFF9FBBFAE5DC3FFC7BCC1FFFFE4F87FFFFF119FF2C21212BFFD023CFDEFE;
defparam prom_inst_24.INIT_RAM_15 = 256'hFFFFFF2B43F5804120959ECCF3F7FFFFFFE69118FEFFFFFFFFFFFFFFC7FFFFED;
defparam prom_inst_24.INIT_RAM_16 = 256'hF932481FFFFFFFFFFFFFFFDFFEEFFBFF8FFFEFF1FEB84F0FA61CBA07FFFF9FDB;
defparam prom_inst_24.INIT_RAM_17 = 256'hFFFDFC2F9F87AFE01F24E0FFFFC5F2FFFFFFE4717E704000F007733EFFFEDFF3;
defparam prom_inst_24.INIT_RAM_18 = 256'hFFFCF66F8E0000DFFFD3FFFF35F9FCFEEFBCEFFFFFFFFFFFFFFFEFEFBEFFCFCE;
defparam prom_inst_24.INIT_RAM_19 = 256'h707BFFFFFFFFFFFFFFFFFBFEFFFBFFFFFFFFD8FFFC2FFC97F9383FFFF3C73FFF;
defparam prom_inst_24.INIT_RAM_1A = 256'h8FF7CDFFCFFF97F0B807FFFCBFDFFFFFFF937FFBC1805FFFFEBFFCFBFBFFF859;
defparam prom_inst_24.INIT_RAM_1B = 256'hF3367F38005FEFFD7FFFFEF7FFDE7E603FEFFFFFFFFFFFFFFEFFFEF7EF26BFFF;
defparam prom_inst_24.INIT_RAM_1C = 256'hFBDFFFFFFFFFFFFFDF8FFC7F47EFFE01BCF81FF2FFCFFC0E01FFFF35D7FFFFFF;
defparam prom_inst_24.INIT_RAM_1D = 256'h1FCFFEFFD1FE4700FFFFCEFDFFFFFFFEB69FEF006F7FFFFE3FBEDFF7E1FBBA82;
defparam prom_inst_24.INIT_RAM_1E = 256'h47F9E1B7FFFFFFDFFFBBFC99DE975030F7FFFFFFFFFFFFFC387F8F90FFFF80F7;
defparam prom_inst_24.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFF87FF81C5FF807F4FF17F6FF43F22007FFFF2067FFFFFFF8C;
defparam prom_inst_24.INIT_RAM_20 = 256'h7FEBF9DFB0001FFFFC1FDFFFFFFFE5F9FF3D5FFFFFFFFFFFFFEFFBFF9F4F1877;
defparam prom_inst_24.INIT_RAM_21 = 256'hE5D6FFFFFFFFDFFFBEDFF887D98BFFFFFFFFFFFFFFFFFF7BFFF0017FE00FF6FE;
defparam prom_inst_24.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFE0005FF003FFFFFE7BF4FBEF000FFFFF9A63FFFFFFF9F67F;
defparam prom_inst_24.INIT_RAM_23 = 256'h7D7ED7E003FFFFE77FFFFFFFFC79DFFC9FBFFFFFFFFBFFFDBFFE21E608FFFFFF;
defparam prom_inst_24.INIT_RAM_24 = 256'h7FFFFFFFF77FFFE7FF85FDE8F03FFFFFFFFFFFFFFFFEFFE00013F800FFE3FD3E;
defparam prom_inst_24.INIT_RAM_25 = 256'hFFFFFFFFFFDFF80071FC003FFDFEBA92BEA5F0007FFFFC759FFFFFFF3C77FF31;
defparam prom_inst_24.INIT_RAM_26 = 256'hEFFC003FFFFF2F43FFFFFF9FEDFFCD1FFFFFFFFFDFFFFFFFFFFE0E134DFFFFFF;
defparam prom_inst_24.INIT_RAM_27 = 256'hFFFFFFFBFFFDFFF79FE7A1FDFFFFFFFFFFFFFFFFFDFC003FEA000BFFFF2F865F;
defparam prom_inst_24.INIT_RAM_28 = 256'hFFFFFFFFFC8C08FE0000FFFD6FF7CFE0FE001FFFFFC7CEFFFFFFEF347FF16F7F;
defparam prom_inst_24.INIT_RAM_29 = 256'h8007FFFFF93EFFFFFFF00ABFFCC3EFFFFFFFE7FFFFFFF5E998082FFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2A = 256'hFFFDFFFFFFA11C6633075FFFFFFFFFFFFFFFFFFF0007FF00000FC790FF9FF93F;
defparam prom_inst_24.INIT_RAM_2B = 256'hFFFFFFDD1B7FD00003C069BFFBFC9F0003FFFFFF33D3FFFFF1FF5FFF37FFFFFF;
defparam prom_inst_24.INIT_RAM_2C = 256'hFFFFFFC7F87FFFF9E727FFCDDFFFFFFFFFDFFFFFFE68FF4468D1FFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2D = 256'hFFFFFFFFF8F6B541EE7FFFFFFFFFFFFFFFFFEFE3FFF80000000007FB7EC68000;
defparam prom_inst_24.INIT_RAM_2E = 256'hFFF7F9BFFF8400000000FEFFF980007FFFFFF91B1FFFF1CDF3FFF15FFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2F = 256'hFFFF3BFBFFF8F959FFFE5DFFFFFFFFFDFFFFFFBE3B6B7879FFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_30 = 256'hFFF9FFFA758281F7FFFFFFFFFFFFFFFFFFFF307F8FF00000001FF78F80003FFF;
defparam prom_inst_24.INIT_RAM_31 = 256'hFE0C0FEFFF0000001BFD8F80000FFFFFFFCB5B7FC75EECFFFF94EFFFFFFFFF3F;
defparam prom_inst_24.INIT_RAM_32 = 256'hF97F704FF5BE7FFFE36FFFFFFFFFE7FFFFFF7D7E07D637FFFFFFFFFFFFFFFFFE;
defparam prom_inst_24.INIT_RAM_33 = 256'hFFBE1F2DFE45FFFFFFFFFFFFFFFFFFBF0187FEFFC0000003AF5FE0003FFFFFFF;
defparam prom_inst_24.INIT_RAM_34 = 256'h7FFE3FF00000003AF9C0000FFFFFFFFE3D0FFF49CD3FFFFCB7FFFFFFFFE9FFFF;
defparam prom_inst_24.INIT_RAM_35 = 256'h6325930B3FFFFF327FFFFFFFF67FFFFFF87F119D97FFFFFFFFFFFFFFFFFFF3C0;
defparam prom_inst_24.INIT_RAM_36 = 256'hFE438EE9BFFFFFFFFFFFFFFFFFFFF83FFFBFFC00000000A8000007FFFFFFFFC9;
defparam prom_inst_24.INIT_RAM_37 = 256'hE07F0000000007000003FFFFFFFFF929F9F58A3FFFFFC64FFEFFFFFA3FFFFF9F;
defparam prom_inst_24.INIT_RAM_38 = 256'hDC963FFFFFF8E9FFFFFFFC17FFFFFF1FBD690BFFFFFFFFFFFFFFFFFFFD5E3FFF;
defparam prom_inst_24.INIT_RAM_39 = 256'h0C423F3FFFFFFFFFFFFFFFFF8B2FFFF20F8000000003F00003FFFFFFFFFF36FE;
defparam prom_inst_24.INIT_RAM_3A = 256'hF000000003FE000FFFFFFFFFFFE1841B167FFFFFFE155FFFFFFF65FFFFFFFFE7;
defparam prom_inst_24.INIT_RAM_3B = 256'h7FFFFBFFC6AE3BFFFFE07FFFFFFFFFC110CFFFFFFFFFFFFFFFFFFFE300FFFFC3;
defparam prom_inst_24.INIT_RAM_3C = 256'h0AFFFFFFFFFFFFFFFFFFF881FFFC70F80000E7DFFFE9DFFFFFFFFFFFFF15B71C;
defparam prom_inst_24.INIT_RAM_3D = 256'h0AFBFFFFFFFFFFFFFFFFFFFFF1FE12FFFFFFFFF8C57DFC7CFF9FFFFFFFE18E50;
defparam prom_inst_24.INIT_RAM_3E = 256'hFF8BFF189F7C1E7EA3FFFFBBF0BE4100D7FFFFFFFFFFFFFFFFFC183FFF8E3E00;
defparam prom_inst_24.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFE0007E80B8F8017FFFFFFFFFFFFFFFFFFFFFFFF80003FFF;

pROM prom_inst_25 (
    .DO({prom_inst_25_dout_w[30:0],prom_inst_25_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_25.READ_MODE = 1'b1;
defparam prom_inst_25.BIT_WIDTH = 1;
defparam prom_inst_25.RESET_MODE = "SYNC";
defparam prom_inst_25.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF07FFFFFBAFFC1AFF7FFBE02FFFFEFFDBE28401F;
defparam prom_inst_25.INIT_RAM_01 = 256'hFFF835FA0E5A003FFFFFBE7C67EC2FFFFFFFFFFFFFFFFFFF80322FF8C78007FF;
defparam prom_inst_25.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFC0067FFE31E003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDE7;
defparam prom_inst_25.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFB8FFFF86597FFC001FFFFEF5FCE5C3866FFF;
defparam prom_inst_25.INIT_RAM_04 = 256'hF86631120003FFFE7CFBA024DEDFFFFFFFFFFFFFFFFFF801CDF5087003FFFFFF;
defparam prom_inst_25.INIT_RAM_05 = 256'hFFFFFFFFFFFE007C960C7C007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCEFF;
defparam prom_inst_25.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFBBFFFF078EE480185FFFFFFFE7C47BE1FFFFFF;
defparam prom_inst_25.INIT_RAM_07 = 256'h1E2D00102BFFF9FFF1F0FFF47FFFFFFFFFFFFFFFFFC01F939D3E00FFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_08 = 256'hFFFFFFFFF801EB7D1F00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF0;
defparam prom_inst_25.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFF7FFFFFF00F1404E057FFF9DFFCE6302FFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_0A = 256'h600844BFFF7FFF1F88487FFFFFFFFFFFFFFFFFFF003D133F803FFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_0B = 256'hFFFFFFD003D87F800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB9FFFFF807;
defparam prom_inst_25.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFF2FEFFFFFFFE03E441C07FFFFFFDFFA140CFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_0D = 256'h0631FFF9B7FFFBE075FFFFFFFFFFFFFFFFFFFC001FFFC01FFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_0E = 256'hFFFFD000FE8007E7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC5EFFFFFFFFFF07C8;
defparam prom_inst_25.INIT_RAM_0F = 256'hFFFFFFFFFFFFFBFF7FFBFFFFFFF87908001FEDEBDC7EF8267FFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_10 = 256'h0BFFFEF1FFFF285FFFFFFFFFFFFFFFFFFFFB00000003C03FFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_11 = 256'hFFE00000008007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF5FD1FFFFBFFFFFF8A3006;
defparam prom_inst_25.INIT_RAM_12 = 256'hFFFFFFFFD9C67FFFFFFFFFFFF9465B80FFFBFFFFA72BFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_13 = 256'hFEEFFFE9E607FFFFFFFFFFFFFFFFFFFFFE0000007C01FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_14 = 256'hF000006FF03FFFFFFFFFFFFFFFFFFFFFFFFFFED6C1FFFFFFFFFFFFFF20C6220F;
defparam prom_inst_25.INIT_RAM_15 = 256'hFFF80A3FFFFFFFFFFFFFFFE4186A04FF9EFF669EF3FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_16 = 256'hFFE7663C9FFFFFFFFFFFFFFFFFFFFFFFA0001FDC0FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_17 = 256'h8016FBE3FFFFFFD17FFFFFFFFFFFFFFCC951FFFFFFFFFFFFFFFFFE821D803FF9;
defparam prom_inst_25.INIT_RAM_18 = 256'h9FFFFFFFFFFFFFFFFFFFD06A1983FBFFFFFBAE1BFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_19 = 256'hFEF6D7FFFFFFFFFFFFFFFFFFFFFFFFF401B788FFFFFFFFFCFFFFFFFFFFFE220D;
defparam prom_inst_25.INIT_RAM_1A = 256'h54733FFFFFBFFFEFFFFFFFFFE015C3FFFFFFFFFFFFFFFFFFFFFA0831027FEFFF;
defparam prom_inst_25.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFF0006C42FFBFFF5D9A6FFFFFFFFFFFFFFFFFFFFFFFFFE03;
defparam prom_inst_25.INIT_RAM_1C = 256'hFEDFFFFFFFFFFFFFFFFFFFFFFFFF81CAB28FFFFFEFFFFFFFFFFFFFE01FFFFFFF;
defparam prom_inst_25.INIT_RAM_1D = 256'hA3FFFFF7FFFFEFFFFFFE0E7FFFFFFFFFFFFFFFFFFFFFFFFFE0090481FEFFFFFF;
defparam prom_inst_25.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFC4C18813FFFFFFCD97DFFFFFFFFFFFFFFFFFFFFFFFFA01F5A;
defparam prom_inst_25.INIT_RAM_1F = 256'h7FFFFFFFFFFFFFFFFFFFFFFFF80B2751FFFFFFFFFFFFFFFFFF05FFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFCA3FFFFFFFFFFFFFFFFF127FFFFFFFF89824007FFFFFEB64B;
defparam prom_inst_25.INIT_RAM_21 = 256'h37FFBFFFFFFFF1348200FFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF817C7DC7F;
defparam prom_inst_25.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFF0372AA3FFFFF9FFFFFFFFFF847FFFFFFFFE0B93007;
defparam prom_inst_25.INIT_RAM_23 = 256'hF7FFFFF7FFE8AFFFFFFFFCAFDF0FFF87F53FFFFFFFFF240D419FFFFFFB7BCFFF;
defparam prom_inst_25.INIT_RAM_24 = 256'hCFFFFFFFFFE4830013FFFFFBFECFFFFFFFFFFFFFFFFFFFFFFFFF83D7E50FFFFF;
defparam prom_inst_25.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFE0CFEA83FFFFFDFFFFFFFFE34FFFFFFFB3E73C03FE1B2C;
defparam prom_inst_25.INIT_RAM_26 = 256'hFFFEFFD28FFFFFFF7F4C1FFFFFFFF8EAFFFFFFFFFD9641007FFFFF7FBFFFFFFF;
defparam prom_inst_25.INIT_RAM_27 = 256'hFFFFFFFFB00480CFFFFFF790FFFFFFFFFFFFFFFFFFFFFFFFF875BD41FFFFFFFF;
defparam prom_inst_25.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFC0E1B20FFFFFFCFFFFEFFD48FFFFFFE3A87FFFFFECF31FF7F;
defparam prom_inst_25.INIT_RAM_29 = 256'h7FC49FFFFFFDEA7FFFFFFBF9DF7184AFFFDFFFF6018801FFFFFF3BBFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_2A = 256'hFFFFFECB21903FFFFDEE7FFFFFFFFFFFFFFFFFFFFFFFFE004EB0FFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_2B = 256'hFFFFFFFFFFFF83EF587FFFFFFE7FFF9FD49FFFFFFCF4FFFFFFFD8EFDDEF107F7;
defparam prom_inst_25.INIT_RAM_2C = 256'h9FFFFFFECBFFFFFFFE43FE7DEC807DCFFFFFD8004067FFFD7BD4FFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_2D = 256'hFFFB008001FFFFFEE7FFFFFFFFFFFFFFFFFFFFFFFFC0F72C1FFFFFFFFFFFEFD4;
defparam prom_inst_25.INIT_RAM_2E = 256'hFFFFFFFFF1B1D60FFFFFFFF3FFFFD49FFFFFFBB3FFFFFFFFACE7F033C0037DFF;
defparam prom_inst_25.INIT_RAM_2F = 256'hFFF587FFFFFFFFE10FFFFF84307DFFFFFF6120583FFFFFEFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_30 = 256'hEC002027FFFF5DFFFFFFFFFFFFFFFFFFFFFFFFF052C907FFFFFFFF7FF7F09FFF;
defparam prom_inst_25.INIT_RAM_31 = 256'hFFFFFC3B7AC3FFFFFFFFDFEFE8CFFFFFF7EFFFFFFFFFE81FFFFFFE6917FFFFFF;
defparam prom_inst_25.INIT_RAM_32 = 256'h8FFFFFFFFFF00FFFFFFFFB21BFFFFFFD804000FFFFF60E7FFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_33 = 256'h900C1FFFFF92DFFFFFFFFFFFFFFFFFFFFFFF0DF961FFFFFFFFF9E3E9C7FFFFEB;
defparam prom_inst_25.INIT_RAM_34 = 256'hFF8C44B0FFFFFFFFFF1BF1E7FFFFEFCFFFFFFFFFF807FFFFFFFF281FFFFFFFB0;
defparam prom_inst_25.INIT_RAM_35 = 256'hFFFFFFFC01FFFFFFFFF685F7FFFFF6001011FFFFBF77FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_36 = 256'h001FFFF9DFFFFFFFFFFFFFFFFFFFFFFFC6FB687FFFFFFFFFFFFBE3FFFFCE1FFF;
defparam prom_inst_25.INIT_RAM_37 = 256'hBDD43FFFFFFFFFFFFDF1FFFFCE9FFFFFFFFFFE01FFFFFFFFFEBC3FFFFFFEC021;
defparam prom_inst_25.INIT_RAM_38 = 256'hFFFF907FFFFFFFFFE907FFFFFFE8440703FFFFFFFFFFFFFFFFFFFFFFFFFFFFE2;
defparam prom_inst_25.INIT_RAM_39 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFF0EDEB0FFFFFFFFFFFFE79FFFFEEBFFFFFFF;
defparam prom_inst_25.INIT_RAM_3A = 256'h87FFFFFFFFFFFF4CFFFFE7BFFFFFFFFFFFF03FFFFFFFFFFEC1FFFFFFFF000A00;
defparam prom_inst_25.INIT_RAM_3B = 256'hF807FFFFFFFFFFDC5FFFFFFFA003800FFFFFFFFFFFFFFFFFFFFFFFFFFFF86625;
defparam prom_inst_25.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC1B7D41FFFFFFFFFFFF867FFFE73FFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_3D = 256'hFFFFFFFFFFC13FFFF63FFFFFFFFFFFFE01FFFFFFFFFFFB07FFFFFFF4220101FF;
defparam prom_inst_25.INIT_RAM_3E = 256'h7FFFFFFFFFFEC0FFFFFFFE8401803FFFF7FFFFFFFFFFFFFFFFFFFFFE05ACB0FF;
defparam prom_inst_25.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFF8F6FD87FFFFFFFFFFFE29FFFF2BFFFFFFFFFFFFFA0;

pROM prom_inst_26 (
    .DO({prom_inst_26_dout_w[30:0],prom_inst_26_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_26.READ_MODE = 1'b1;
defparam prom_inst_26.BIT_WIDTH = 1;
defparam prom_inst_26.RESET_MODE = "SYNC";
defparam prom_inst_26.INIT_RAM_00 = 256'hFFFFFFF14FFFFB5FFFFFFFFFFFFFECBFFFFFFFFFFFD03FFFFFFFD000230FFFFF;
defparam prom_inst_26.INIT_RAM_01 = 256'hFFFFFFFFFBC7FFFFFFFA0A80C0FFFFFFFFFFFFFFFFFFFFFFFFFF83A1D41FFFFF;
defparam prom_inst_26.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFE0F8EB0FFFFFFFFFFFF8A3FFF88FFFFFFFFFFFFFF20FFF;
defparam prom_inst_26.INIT_RAM_03 = 256'hFFFC91FFFE57FFFFFFFFFFFFFCC3FFFFFFFFFFFE607FFFFFFF4002C19FFFFFFF;
defparam prom_inst_26.INIT_RAM_04 = 256'hFFFFFFDC1FFFFFFFE8000127FFFFFFFFFFFFFFFFFFFFFFFFE0DD7583FFFFFFFF;
defparam prom_inst_26.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFF07C5741FFFFFFFFFFFE14FFFE6BFFFFFFFFFFFFFF7AFFFFFF;
defparam prom_inst_26.INIT_RAM_06 = 256'h823FFF14FFFFFFFFFFFFFFDE3FFFFFFFFFFFF7DFFFFFFFFD058020FFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_07 = 256'hFFFEB1FFFFFFFFA080E04FFFFFFFFFFFFFFFFFFFFFFFFC0ADEB03FFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_08 = 256'hFFFFFFFFFFF81E66583FFFFFFFFFFFC51FFF8C7FFFFFFFFFFFFFF983FFFFFFFF;
defparam prom_inst_26.INIT_RAM_09 = 256'hFFC41FFFFFFFFFFFFFFE60FFFFFFFFFFFFDC3FFFFFFFF0013813FFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0A = 256'hF787FFFFFFFE0060187FFFFFFFFFFFFFFFFFFFFFFC0CE3A40FFFFFFFFFFFE09F;
defparam prom_inst_26.INIT_RAM_0B = 256'hFFFFFFFC03D4EB03FFFFFFFFFFF04FFFE34FFFFFFFFFFFFFFF9A3FFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0C = 256'hA3FFFFFFFFFFFFFFF7FFFFFFFFFFFFFEF1FFFFFFFFC0003007FFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0D = 256'h7FFFFFFFF8001E0CFFFFFFFFFFFFFFFFFFFFFC01F5F580FFFFFFFFFFF973FFF0;
defparam prom_inst_26.INIT_RAM_0E = 256'hFFFE007432407FFFFFFFFFFC29FFF871FFFFFFFFFFFFFFFC60FFFFFFFFFFFFBC;
defparam prom_inst_26.INIT_RAM_0F = 256'hFFFFFFFFFFFFFF9C7FFFFFFFFFFFF40FFFFFFFFF0038080FFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_10 = 256'hFFFFFFE0640801FFFFFFFFFFFFFFFFFFFE003F7AB03FFFFFFFFFFE047FFC707F;
defparam prom_inst_26.INIT_RAM_11 = 256'h00DCBF580FFFFFFFFFFF823FFE123FFFFFFFFFFFFFFFEFCFFFFFFFFFFFFC13FF;
defparam prom_inst_26.INIT_RAM_12 = 256'hFFFFFFFFFFFDF9FFFFFFFFFFFF40FFFFFFFFFC0004067FFFFFFFFFFFFFFFFFFE;
defparam prom_inst_26.INIT_RAM_13 = 256'hFFFF8008C20FFFFFFFFFFFFFFFFFFE03E4E32403FFFFFFFFFFC28FFF0D0FFFFF;
defparam prom_inst_26.INIT_RAM_14 = 256'h83FB00FFFFFFFFFFE347FF86C3FFFFF7FFFFFFFFFF263FFFFFFFFFFFC07FFFFF;
defparam prom_inst_26.INIT_RAM_15 = 256'hFFFFFFFFF3FFFFFFFFFFFFE01FFFFFFFFFF01904C0FFFFFFFFFFFFFFFFFBBF33;
defparam prom_inst_26.INIT_RAM_16 = 256'hFE6402808FFFFFFFFFFFFFFFFF8FFD3855C07FFFFFFFFFF963FFE3A1FFFFFFFF;
defparam prom_inst_26.INIT_RAM_17 = 256'h701FFFFFFFFFFE28FFF010FFFFFFFFFFFFFFFFFEFF7FFFFFFFFFF107FFFFFFFF;
defparam prom_inst_26.INIT_RAM_18 = 256'hFFFFFF9FDFFFFFFFFFFDC1FFFFFFFFFFD0041087FFFFFFFFFFFFFFFA07AF77F2;
defparam prom_inst_26.INIT_RAM_19 = 256'h8DC0607FFFFFFFFFFFFFFB02C6ED9E9807FFFFFFFFFF243FF8683FFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_1A = 256'hFFFFFFFFFF903FFE365FFFFFFFFFFFFFFFFFF270FFFFFFFFFE00FFFFFFFFFFFA;
defparam prom_inst_26.INIT_RAM_1B = 256'hFFFF3F9FFFFFFFFF807FFFFFFFFFFF5201604FFFFFFFFFFFFFFC780746256E00;
defparam prom_inst_26.INIT_RAM_1C = 256'h2001FFFFFFFFFFFFFF6073EE56D3C01FFFFFFFFFC68FFE0B07FFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_1D = 256'hFFFFFFF203FF0281FFFFFFFFFFFFFFFFFFEBF7FFFFFFFF8C1FFFFFFFFFFFEE01;
defparam prom_inst_26.INIT_RAM_1E = 256'hF9ACBFFFFFFF0027FFFFFFFFFFFDC040283FFFFFFFFFFFFF403BED331A7807FF;
defparam prom_inst_26.INIT_RAM_1F = 256'h07FFFFFFFFFFFF100FF9C780DE00FFFFFFFFF891FFC1617FFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_20 = 256'hFFFC48FFE0505FFFFFFFFFFFFFFFFFFF17FEFFFFFEFE03FFFFFFFFFFFFA8C034;
defparam prom_inst_26.INIT_RAM_21 = 256'hFFDEFFF97321FFFFFFFFFFFFF5001608FFFFFFFFFFFF8023F2F6A019C01FFFFF;
defparam prom_inst_26.INIT_RAM_22 = 256'hFFFFFFFFFFC211FD94F006780FFFFFFFFF123FF02C0FFFFFFFFFFFFFFFFFFFE2;
defparam prom_inst_26.INIT_RAM_23 = 256'hC81FF81A03FFFFFFFFFFFFFFFFFFFE47FFDEB9FE79FFFFFFFFFFFFFCE039080F;
defparam prom_inst_26.INIT_RAM_24 = 256'hFFFFE7FCFFFFFFFFFFFFFFD41E11A1FFFFFFFFFFE08476FCAC00E603FFFFFFFF;
defparam prom_inst_26.INIT_RAM_25 = 256'hFFFFFFF8687F7E27002DC0FFFFFFFFE0C7FE0D83FFFFFFFFFFFFFFFFFFFF86DD;
defparam prom_inst_26.INIT_RAM_26 = 256'hFF03C03FFFFFFFFFFFFFFFFFF6B85A1DDE7DF87FFFFFFFFFFFFFFA8008067FFF;
defparam prom_inst_26.INIT_RAM_27 = 256'hFFF8FFFFFFFFFFFFFFFE501C4687FFFFFFFFFC1A7FBFB58004303FFFFFFFF803;
defparam prom_inst_26.INIT_RAM_28 = 256'hFFFE0E3FDFA898632C17FFFFFFFE18FF80E01FFFFFFFFFFFFFF6F7281A0C327F;
defparam prom_inst_26.INIT_RAM_29 = 256'h3807FFFFFFFFFFFFD0400204B80C3F7CE0FFFFFFFFFFFFFFFFCE150021FFFFFF;
defparam prom_inst_26.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFD4607007FFFFFFFFF03EF6FEB7C00DB01FFFFFFFF107F80;
defparam prom_inst_26.INIT_RAM_2B = 256'h81FFD7F5CF002C407FFFFFFFCB1FF01603FFFFFFFFFFFFE0000D00308008E773;
defparam prom_inst_26.INIT_RAM_2C = 256'h7FEFFFFFFFFE000000400355000007FFFFFFFFFFFFFFFFFF08009007FFFFFFFF;
defparam prom_inst_26.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFE500DC01FFFFFFFFF0E7F57FA3000EB01FFFFFFFF08BF00500;
defparam prom_inst_26.INIT_RAM_2E = 256'h7D3E0FC005EC03FFFFFFFC03FC03C017FF7FFFFFFF000019200011B200FFFFFF;
defparam prom_inst_26.INIT_RAM_2F = 256'hDFFFFFDA00001C00000804E7FFFFFFFFFFFFFFFFFFFFFCA470007FFFFFFFF878;
defparam prom_inst_26.INIT_RAM_30 = 256'hFFFFFFFFFFFF9C40001FFFFFFFFC105F794FE001CA00FFFFFFFE58E400B001BF;
defparam prom_inst_26.INIT_RAM_31 = 256'h2C7000F980DFFFFFFF0076806C007FFFFFFFF680001CA10000945BFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_32 = 256'hFFC380001E7190000522FFFFFFFFFFFFFFFFFFFFFFF1800007FFFFFFFC26BFCA;
defparam prom_inst_26.INIT_RAM_33 = 256'hFFFFFFFFFE700001FFFFFFFF4127FDA1780059600FFFFFFFE01D000E001EFFBF;
defparam prom_inst_26.INIT_RAM_34 = 256'h006FB001FFFFFFD844C0038003FEFFFFFE00000F193D14004E07FFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_35 = 256'h00000F84FFD2803407FFFFFFFFFFFFFFFFFFFFFFE300007FFFFFFA6029CF3FF4;
defparam prom_inst_26.INIT_RAM_36 = 256'hFFFFFFFD00003FFFFFFE685487D86500268C00FFFFFFFC700001E000FFFFFFF6;
defparam prom_inst_26.INIT_RAM_37 = 256'h56003FFFFFFC20000058000FFFFFFF800007DB77F52802407FFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_38 = 256'h01E3DBFF9E80EA0FFFFFFFFFFFFFFFFFFFFFFF88005FFFFFFFB0448921100077;
defparam prom_inst_26.INIT_RAM_39 = 256'hFFFFF9F827FFFFFF34280008A30001EB000FFFFFFFA2000016000BFFFF9EB800;
defparam prom_inst_26.INIT_RAM_3A = 256'h07BFFFFFC08080050011FFFFF7D00001F5EDFFC1F80C81FFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3B = 256'h26FFFF6F81C80FFFFFFFFFFFFFFFFFFFFFFF87DFFFFFFF3F1F1E20008009D580;
defparam prom_inst_26.INIT_RAM_3C = 256'hFFFF1FFFFFFFCFFE2720150005EAC001FFFFFF8160000340043BFFEFBA0000F8;
defparam prom_inst_26.INIT_RAM_3D = 256'hFFF7A008000078010FB7FB8E00007D73FFFFF7D82881FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3E = 256'hFBFF5D83887FFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFCFCFF1E112A0017160007F;
defparam prom_inst_26.INIT_RAM_3F = 256'hFFFFFFFFE7F3BCFE05C001BCB00003FFFFFE1400001C00023FED8000007E0FDF;

pROM prom_inst_27 (
    .DO({prom_inst_27_dout_w[30:0],prom_inst_27_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_27.READ_MODE = 1'b1;
defparam prom_inst_27.BIT_WIDTH = 1;
defparam prom_inst_27.RESET_MODE = "SYNC";
defparam prom_inst_27.INIT_RAM_00 = 256'h0000000931EDFFFFFFFFFFFFFFFFBFFFFFFF679FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_01 = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB800000;
defparam prom_inst_27.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFF600000000000000403F7EFFFF767FFDFF87DBFFFF;
defparam prom_inst_27.INIT_RAM_03 = 256'h000021597FFFFFFFFFFFFCFFBA7FFFFFDC6DBFFFFFFFFFFFFFFFFFFFFFFFEFFF;
defparam prom_inst_27.INIT_RAM_04 = 256'hE7DDD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1000007800;
defparam prom_inst_27.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFEC00000700000000001397DFFF9FFFFFFC819F61D8007;
defparam prom_inst_27.INIT_RAM_06 = 256'h0000184EF7FE79FFFF300210006001999A76FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_07 = 256'hE0FCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFED0000020000000;
defparam prom_inst_27.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFBE400000300060000000021B79DFFFFF4C0208100108032B43;
defparam prom_inst_27.INIT_RAM_09 = 256'h0100637FB41E8600000040400B664A2D02CFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_0A = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB2080000580004000000;
defparam prom_inst_27.INIT_RAM_0B = 256'hFFFFFFFFFFEF420000100001C00000005818FFE807A0800008205002C86A8860;
defparam prom_inst_27.INIT_RAM_0C = 256'h01FF8696003008200000001049C0027FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7400000E00007F00000000;
defparam prom_inst_27.INIT_RAM_0E = 256'hFFFFFFFFFB000007E000F860000108007FE020800C0100000000001A800037FF;
defparam prom_inst_27.INIT_RAM_0F = 256'hFE068000000200000000184E081FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF3400009FE00FE0E000000241F;
defparam prom_inst_27.INIT_RAM_11 = 256'hFFFFFD0080041FF03C00F000100539F786440C000000002000038AEF0DFCFFFF;
defparam prom_inst_27.INIT_RAM_12 = 256'h910300000000000000622DC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBB40400E01FE7F000EA04100CFFBE1;
defparam prom_inst_27.INIT_RAM_14 = 256'hFFA4000C001FFF00006007F9FE7FDB837000000000001080009D1C73FFFFFFFF;
defparam prom_inst_27.INIT_RAM_15 = 256'h10000C000008000001844F5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000F0001F700000D3FF7DFFFFDF962;
defparam prom_inst_27.INIT_RAM_17 = 256'h800200003AE0001F5FFFFFFFFEEFF88000F000000000000042EC5FEFFFEFEFFF;
defparam prom_inst_27.INIT_RAM_18 = 256'h0240018100000000F8FFFDFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_27.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB680580002E3E000FC1FFFFFFEFFF7A0000;
defparam prom_inst_27.INIT_RAM_1A = 256'hF8001F8FE00F801FFFEFFFFFE6C00000000068400000602233FFFFBFFFBFFFFF;
defparam prom_inst_27.INIT_RAM_1B = 256'h0000800000003D3FDAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC400;
defparam prom_inst_27.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFBF1275F0017C0FE03E001FDFFFFFFFE60000000;
defparam prom_inst_27.INIT_RAM_1D = 256'h0FE01FF7C0001BFFFFFFFFE00000000101010000000B0EFFCFFFFFFF7FFFFFFF;
defparam prom_inst_27.INIT_RAM_1E = 256'hC0A0000002C3FFDFDFEFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEB60C3F0;
defparam prom_inst_27.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFBF1C07F0FC000FFF00003FFFFFFFFF8000000FF01;
defparam prom_inst_27.INIT_RAM_20 = 256'h0007F80000FFFFFFFF7618000BFCD1400055002020FFAFFFF7FFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_21 = 256'h0100004F97DFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFCC007F3F0;
defparam prom_inst_27.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFBFE0007FE00003EE0001F7FFFFFFF4800005F8018200;
defparam prom_inst_27.INIT_RAM_23 = 256'hF7E00077FFFFFFF6400001F8873C000025010307FBFFFBFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_24 = 256'h40016FDFDBFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBC00007D00003;
defparam prom_inst_27.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFF3F00003F78001F8FF00F8FFFFFFFF400003F0112D800000;
defparam prom_inst_27.INIT_RAM_26 = 256'hF0383FFFFFFE480003F02215E00000100269F7F9FBFDFFEFFFF7FFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_27 = 256'h000FFDFFF77B3FE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCDC0002FEF801FE0F;
defparam prom_inst_27.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFEFC001FDBF81BF00FFFD0FFFFFFFF00020700EB03E00000400;
defparam prom_inst_27.INIT_RAM_29 = 256'h03FFFFFFFC80003818640EE0000000000EDFFFBCFCD97FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2A = 256'h87FFFF3F33DFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7C017A07FE7E000FFF;
defparam prom_inst_27.INIT_RAM_2B = 256'hFFFFFFFFFFFF1FC1FC007FDF0000FE80FFFFFFFD20001E0802300E0000000003;
defparam prom_inst_27.INIT_RAM_2C = 256'hFFFFFFA00007C0C0400190000000001EEFFE7FF7B9FFFBFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2D = 256'hF3FFFFBFEEDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7CBE0007FF00001F003F;
defparam prom_inst_27.INIT_RAM_2E = 256'hFFFFFFFFFFF7FE0000FFF0000F100FFFFFFFD60043F82080007C00000000003C;
defparam prom_inst_27.INIT_RAM_2F = 256'hFFE60200FF0480000F00000000000C3E7FDBDDFBF1FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_30 = 256'hB7FEFFEEFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F00007FFC0007B403FFFF;
defparam prom_inst_27.INIT_RAM_31 = 256'hFFFFFFEFFF80003FFF4005EC00FFFFFFFD40003FE10000F7F00000000000BF3F;
defparam prom_inst_27.INIT_RAM_32 = 256'hD0203FFCE001E4FD00005880001FCFFFE6BEFBDFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_33 = 256'h9EFE7FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFBFE78000FD7FC03C100DFFFFFFF;
defparam prom_inst_27.INIT_RAM_34 = 256'hFFFF7F9F802FF1FF42E04007FFFFFFF800017FB003FC1F80001DEA01004DFFFB;
defparam prom_inst_27.INIT_RAM_35 = 256'h0017F0031401F80008001080C3EEF597FCFFFEFFFBFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_36 = 256'h6167FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE5F80DE00FF1E00025FFFFFFFFC0;
defparam prom_inst_27.INIT_RAM_37 = 256'hFFF8DF87F801FFF00122FFFFFFFFF00047FC8319D83E000580062433F8BFE3FE;
defparam prom_inst_27.INIT_RAM_38 = 256'hFFB110702FA00026020026DCFDFBF7FCDF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_39 = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF7E1FFEF00007FC00201FFFFFFDDC284F;
defparam prom_inst_27.INIT_RAM_3A = 256'hCFFFFC2001F400400FFFFFFFFF5D73FFF6206360F80000002001A37FFF4FFFAF;
defparam prom_inst_27.INIT_RAM_3B = 256'h8C60801F000000002037FFEFE77FA7E76B3FFFFFFFFFFFFFFFFFFFFFFFFFFFC7;
defparam prom_inst_27.INIT_RAM_3C = 256'hFDFFFFFFFFFFFFFFFFFFFFFFFFFFF973FFFC00405E001081FFFFFFFFFFDDFFFE;
defparam prom_inst_27.INIT_RAM_3D = 256'hDFF0003C800400FFFFFFFFFFFFFFFFE6818CC3F00000000058CCFFFE19E76E1B;
defparam prom_inst_27.INIT_RAM_3E = 256'h82803C0000000026333FFF9E79D9E3FF7FFFFFFFFFFFFFFFFFFFFFFFFFFE963F;
defparam prom_inst_27.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF91FFAF8002F0003000FFFFFFFFFFFFFFFFE50;

pROM prom_inst_28 (
    .DO({prom_inst_28_dout_w[30:0],prom_inst_28_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_28.READ_MODE = 1'b1;
defparam prom_inst_28.BIT_WIDTH = 1;
defparam prom_inst_28.RESET_MODE = "SYNC";
defparam prom_inst_28.INIT_RAM_00 = 256'hC01E0103000BFFFFFFFFFFFBFFFFCA011347C00000800B40FEF5F87E4423314F;
defparam prom_inst_28.INIT_RAM_01 = 256'h00F00000000037FEFFBFE7E3F93D77FFFFFFFFFFFFFFFFFFFFFFFFFFEB83FF0F;
defparam prom_inst_28.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFBE1FF8CFC3F42401403FFFFFFFFFEF8B8FFFD4208;
defparam prom_inst_28.INIT_RAM_03 = 256'hC04194017FFFFFFFFF12763FFF280C0D3F0000000004FF9FEB79F167BEFF6FFF;
defparam prom_inst_28.INIT_RAM_04 = 256'hE0000000848EBDFFFFF03877DFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FF1CFCB;
defparam prom_inst_28.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFC0FC7CFFA03089003FFFFFFFFF8618767FF4040407;
defparam prom_inst_28.INIT_RAM_06 = 256'h4440CFFFFFFFFE60800C0FFEC01812FE00000002236F779F7B873FF9FFFFFFFF;
defparam prom_inst_28.INIT_RAM_07 = 256'h000000015FFFDEFE40817EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8BD0FCFE00C;
defparam prom_inst_28.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFF37E3FCF00104107AFFFFFFFF1C0C2019BFC810541FE0;
defparam prom_inst_28.INIT_RAM_09 = 256'h0BBFFFFFBF201B06025BF9006C09FC000000003FFDFFFFF967FFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0A = 256'h000C3FFFFFFFE6187FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF867AFFD0008204;
defparam prom_inst_28.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFF1F3ED1FF100220121EFFFFFFF802701780F7F2018D83F8000;
defparam prom_inst_28.INIT_RAM_0C = 256'hFFFFFFF33C3F0F819FE4002007F02000002DFFFFF8E011F978DEFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0D = 256'h13FFDF9E7F1AED1FFF7FFFFFFFFFFFFFFFFFFFF7FFFFFC1E7FCFFC001480439B;
defparam prom_inst_28.INIT_RAM_0E = 256'hFFFF7FFFFFFFE10FEEFF800820114EFFFFFFF454FFFC4E02FC800130FF400100;
defparam prom_inst_28.INIT_RAM_0F = 256'hFFF800FFFFE341DF9020A00FF00000009FF7FFDF9F78A7EFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_10 = 256'hDFFFFDE7A0F8DDFFFFFFFFFFFFFFFFEFFFDFBF37FFFE23FF5FE20C801C23BFFF;
defparam prom_inst_28.INIT_RAM_11 = 256'hFFEFBFFFFBE0FFDFFA86180420DFFFFFFF757FFFFF28EFF200C0D1FFFB0003DF;
defparam prom_inst_28.INIT_RAM_12 = 256'h1DBFFFFFF202FE4080007FFE4200FFF4FFFEFFF90F375FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_13 = 256'hFFFFF3847F7DFFFFFFFFFFFFFFFEFFFFFBFFFFFEFC3FE1DE8042806867FFFFFF;
defparam prom_inst_28.INIT_RAM_14 = 256'hFFF7FFDF8BFDD9E301A34A3BFFFFFF901FFFFFFE601FC8012127FFD023CFDEFE;
defparam prom_inst_28.INIT_RAM_15 = 256'hFFFFFFC43DF900476058BECCF3F7FFFFFFE69118FEFFFFFFFFFFFFFFB7FFBFBD;
defparam prom_inst_28.INIT_RAM_16 = 256'hF932481FFFFFFFFFFFFFFFDF7FEFFBFFFDFFFFF87E3B80106122C9FFFFFFEC37;
defparam prom_inst_28.INIT_RAM_17 = 256'hFFFFFC17AFB8101110B91FFFFFFA09FFFFFFF94EFFA040C08FF9733EFFFEDFF3;
defparam prom_inst_28.INIT_RAM_18 = 256'hFFFF281FF4018020002BFFFF35F9FCFEEFBCEFFFFFFFFFFFFFFFFFEFBFFEDFDE;
defparam prom_inst_28.INIT_RAM_19 = 256'h707BFFFFFFFFFFFFFFFBFFFFFFBBF6FFFFBFDF31FBC800181EC7FFFFFD38FFFF;
defparam prom_inst_28.INIT_RAM_1A = 256'hF7E7F0FFF400C80047FFFFFF403FFFFFFFE603FC8180A060017FFCFBFBFFF859;
defparam prom_inst_28.INIT_RAM_1B = 256'hFDC9FFD00020080387FFFEF7FFDE7E603FEFFFFFFFFFFFFFFFFFFEFDCFB3BFFF;
defparam prom_inst_28.INIT_RAM_1C = 256'hFBDFFFFFFFFFFFFFDFFBFFFFFFFFFFFE7CFBDFF500140171FFFFFFD80FFFFFFF;
defparam prom_inst_28.INIT_RAM_1D = 256'hBFB7FD003001B8FFFFFFF503FFFFFFFF213FF20050900001FFBEDFF7E1FBBA82;
defparam prom_inst_28.INIT_RAM_1E = 256'h1FFE41482000002FFFBBFC99DE975030F7FFFFFFFFFFFFFFBFD7FFFFFFFFFF03;
defparam prom_inst_28.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFF7FFFFFFFDFFFF800FF67F001040DDFFFFFFFC99FFFFFFFFE8;
defparam prom_inst_28.INIT_RAM_20 = 256'h8FF000506FFFFFFFFFA03FFFFFFFFB03FFC9A000000000FFFFEFFBFF9F4F1877;
defparam prom_inst_28.INIT_RAM_21 = 256'hF969000000003FFFBEDFF887D98BFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFF006FE;
defparam prom_inst_28.INIT_RAM_22 = 256'hFFFFFFFFFFFFEFFFFFFFDFFFFC007FC0780C9820FFFFFFFFEC17FFFFFFFE88FF;
defparam prom_inst_28.INIT_RAM_23 = 256'hA402201FFFFFFFFA81FFFFFFFF863FFF264000000003FFFDBFFE21E608FFFFFF;
defparam prom_inst_28.INIT_RAM_24 = 256'h8000000008FFFFE7FF85FDE8F03FFFFFFFFFFFFFFFFEFFFFFFFFFFFF0013F9CF;
defparam prom_inst_28.INIT_RAM_25 = 256'hFFFFFFFFFFDFFFFF8CFFFFC002FD3CAC409A0FFFFFFFFF427FFFFFFFC01FFFC4;
defparam prom_inst_28.INIT_RAM_26 = 256'h6C03FFFFFFFFC81FFFFFFFE01BFFF1A0000000001FFFFFFFFFFE0E134DFFFFFF;
defparam prom_inst_28.INIT_RAM_27 = 256'h00000007FFFDFFF79FE7A1FDFFFFFFFFFFFFFFFFFDFFFFC05FFFF4000F4FC800;
defparam prom_inst_28.INIT_RAM_28 = 256'hFFFFFFFFFD7FF003FFFF0002E7F0101101FFFFFFFFFB00FFFFFFF0C9FFFE6080;
defparam prom_inst_28.INIT_RAM_29 = 256'h7FFFFFFFFE611FFFFFFD107FFF0C1000000018FFFFFFF5E998082FFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2A = 256'h00023FFFFFA11C6633075FFFFFFFFFFFFFFFFFFEFFF800FFFFF0386EFF6004C0;
defparam prom_inst_28.INIT_RAM_2B = 256'hFFFFFFE3FC002FFFFC3F963FF00360FFFFFFFFFFD8E7FFFFFF003FFFC5000000;
defparam prom_inst_28.INIT_RAM_2C = 256'hFFFFFFFA01FFFFFE18DFFFF1E00000000027FFFFFE68FF4468D1FFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2D = 256'h01FFFFFFF8F6B541EE7FFFFFFFFFFFFFFFFFD01C0003FFFFFFFFFFF881B97FFF;
defparam prom_inst_28.INIT_RAM_2E = 256'hFFF80600017BFFFFFFFEFE20C67FFFFFFFFFFE60FFFFFE022FFFFE5000000000;
defparam prom_inst_28.INIT_RAM_2F = 256'hFFFFD40FFFFF00B7FFFF9600000000027FFFFFBE3B6B7879FFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_30 = 256'hFFF9FFFA758281F7FFFFFFFFFFFFFFFFFE00CF80400FFFFFFFFFC8107FFFFFFF;
defparam prom_inst_28.INIT_RAM_31 = 256'h01F3F01800FFFFFFE5F8607FFFFFFFFFFFF2BCFFFC801BFFFFE61000000000DF;
defparam prom_inst_28.INIT_RAM_32 = 256'hFE426BB00075FFFFFDA0000000001FFFFFFF7D7E07D637FFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_33 = 256'hFFBE1F2DFE45FFFFFFFFFFFFFFFFFFE0FE7802003FFFFFFC5C301FFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_34 = 256'h8001800FFFFFFFC50E3FFFFFFFFFFFFFDA8000303CFFFFFF240000000017FFFF;
defparam prom_inst_28.INIT_RAM_35 = 256'h89C200E8FFFFFFC4800000000AFFFFFFF87F119D97FFFFFFFFFFFFFFFFFFFC3F;
defparam prom_inst_28.INIT_RAM_36 = 256'hFE438EE9BFFFFFFFFFFFFFFFFFFD07C0005003FFFFFFFF43FFFFFFFFFFFFFFF3;
defparam prom_inst_28.INIT_RAM_37 = 256'h1800FFFFFFFFFFFFFFFFFFFFFFFFFE4A000079FFFFFFF89001000004BFFFFF9F;
defparam prom_inst_28.INIT_RAM_38 = 256'h0751FFFFFFFF32000000036FFFFFFF1FBD690BFFFFFFFFFFFFFFFFFFFFA1C000;
defparam prom_inst_28.INIT_RAM_39 = 256'h0C423F3FFFFFFFFFFFFFFFFFECF0000E007FFFFFFFFFFFFFFFFFFFFFFFFFC701;
defparam prom_inst_28.INIT_RAM_3A = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFE2B26F1FFFFFFFFE640000000FBFFFFFFFFE7;
defparam prom_inst_28.INIT_RAM_3B = 256'hFFFFFBFFF8C80000001FFFFFFFFFFFC110CFFFFFFFFFFFFFFFFFFFFDFF0001C0;
defparam prom_inst_28.INIT_RAM_3C = 256'h0AFFFFFFFFFFFFFFFFFFFFBE0003F007FFFFFFFFFFFFFFFFFFFFFFFFFFE678D3;
defparam prom_inst_28.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0011FFFFFFFFFF09000380007FFFFFFFE18E50;
defparam prom_inst_28.INIT_RAM_3E = 256'hFF8BFFE12083E002AFFFFFBBF0BE4100D7FFFFFFFFFFFFFFFFFFFFC000FE01FF;
defparam prom_inst_28.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFCF80BDF807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF;

pROM prom_inst_29 (
    .DO({prom_inst_29_dout_w[30:0],prom_inst_29_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_29.READ_MODE = 1'b1;
defparam prom_inst_29.BIT_WIDTH = 1;
defparam prom_inst_29.RESET_MODE = "SYNC";
defparam prom_inst_29.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBAFFFE3400000203FFFFEFFDBE28401F;
defparam prom_inst_29.INIT_RAM_01 = 256'hFFFFC645F006003FFFFFBE7C67EC2FFFFFFFFFFFFFFFFFFFFFCF9FFFC07FFFFF;
defparam prom_inst_29.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFF8DFFCF01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDE7;
defparam prom_inst_29.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFB8FFFFF86180040007FFFEF5FCE5C3866FFF;
defparam prom_inst_29.INIT_RAM_04 = 256'hFF87C2220008FFFE7CFBA024DEDFFFFFFFFFFFFFFFFFFFFE0DFF380FFFFFFFFF;
defparam prom_inst_29.INIT_RAM_05 = 256'hFFFFFFFFFFFFFF80EF9403FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCEFF;
defparam prom_inst_29.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFBBFFFFF80F4080103FFFFFFFE7C47BE1FFFFFF;
defparam prom_inst_29.INIT_RAM_07 = 256'hE038802807FFF9FFF1F0FFF47FFFFFFFFFFFFFFFFFFFE0194B01FFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_08 = 256'hFFFFFFFFFFFE03FB00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFF;
defparam prom_inst_29.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFF03C06804FFFF9DFFCE6302FFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_0A = 256'h4040081FFF7FFF1F88487FFFFFFFFFFFFFFFFFFFFFC00F007FFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_0B = 256'hFFFFFFFFFC18007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB9FFFFFFF8;
defparam prom_inst_29.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFEFEFFFFFFFFFCA000403FFFFFFDFFA140CFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_0D = 256'h35107FF9B7FFFBE075FFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_0E = 256'hFFFFFFFF017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBA0FFFFFFFFFFF940;
defparam prom_inst_29.INIT_RAM_0F = 256'hFFFFFFFFFFFFFC00BFFBFFFFFFFFA82C060FEDEBDC7EF8267FFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_10 = 256'h09FFFEF1FFFF285FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC83BFFFFBFFFFFFF00002;
defparam prom_inst_29.INIT_RAM_12 = 256'hFFFFFFFFF0EDFFFFFFFFFFFFFE000A883FFBFFFFA72BFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_13 = 256'hFEEFFFE9E607FFFFFFFFFFFFFFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_14 = 256'hFFFFFF102FFFFFFFFFFFFFFFFFFFFFFFFFFFFF023FFFFFFFFFFFFFFFC8360107;
defparam prom_inst_29.INIT_RAM_15 = 256'hFFF419FFFFFFFFFFFFFFFFF9000805FF9EFF669EF3FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_16 = 256'hFFE7663C9FFFFFFFFFFFFFFFFFFFFFFFFFFFC445FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_17 = 256'hFFE73E9FFFFFFFE0FFFFFFFFFFFFFFFF80CFFFFFFFFFFFFFFFFFFF2015041FF9;
defparam prom_inst_29.INIT_RAM_18 = 256'h7FFFFFFFFFFFFFFFFFFFE41A0887FBFFFFFBAE1BFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_19 = 256'hFEF6D7FFFFFFFFFFFFFFFFFFFFFFFFFFF7D7E7FFFFFFFFFCFFFFFFFFFFFF401C;
defparam prom_inst_29.INIT_RAM_1A = 256'hCC88FFFFFFFFFFE7FFFFFFFFF80C3FFFFFFFFFFFFFFFFFFFFFFC800402FFEFFF;
defparam prom_inst_29.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFD00A861FFBFFF5D9A6FFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_29.INIT_RAM_1C = 256'hFEDFFFFFFFFFFFFFFFFFFFFFFFFFFF17667FFFFFFFFFFF7FFFFFFF817FFFFFFF;
defparam prom_inst_29.INIT_RAM_1D = 256'h9FFFFFFFFFFFFFFFFFFF85FFFFFFFFFFFFFFFFFFFFFFFFFFFA010403FEFFFFFF;
defparam prom_inst_29.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFF0002017FFFFFFCD97DFFFFFFFFFFFFFFFFFFFFFFFFFFF97D;
defparam prom_inst_29.INIT_RAM_1F = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFEB8CFFFFFFFFFFFFDFFFFFC13FFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_20 = 256'hFFFF7FFFFFFFFFF86FFFFFFFFFFFFFFFFFFDB9FFFFFFFFE004630FFFFFFEB64B;
defparam prom_inst_29.INIT_RAM_21 = 256'h38007FFFFFFFFC008241FFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE43C33FF;
defparam prom_inst_29.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFF9AE59FFFFFFDFFFFFFFFFF0DFFFFFFFFFFEC70FF8;
defparam prom_inst_29.INIT_RAM_23 = 256'hF7FFFFFFFFF19FFFFFFFFF703FF0007E0CDFFFFFFFFF800001BFFFFFFB7BCFFF;
defparam prom_inst_29.INIT_RAM_24 = 256'h3FFFFFFFFFF0003187FFFFFBFECFFFFFFFFFFFFFFFFFFFFFFFFFFC2F1CFFFFFF;
defparam prom_inst_29.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFB9E7FFFFFFFFFFFFBFFE13FFFFFFFEC1303FC00003C;
defparam prom_inst_29.INIT_RAM_26 = 256'hFFFFFFE27FFFFFFFA2C3FFFFFC00021DFFFFFFFFFE044120FFFFFF7FBFFFFFFF;
defparam prom_inst_29.INIT_RAM_27 = 256'hFFFFFFFFC00020DFFFFFF790FFFFFFFFFFFFFFFFFFFFFFFFFF8BCB3FFFFFFF7F;
defparam prom_inst_29.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFF1E11FFFFFFFEFFFFE7FE07FFFFFFF4E7FFFFFFF30CE009F;
defparam prom_inst_29.INIT_RAM_29 = 256'h3FE07FFFFFFE89FFFFFFFC06208E7B6FFFDFFFF80018C3FFFFFF3BBFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2A = 256'hFFFFFF0221807FFFFDEE7FFFFFFFFFFFFFFFFFFFFFFFFFF7B18FFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2B = 256'hFFFFFFFFFFFFFCF8C7FFFFFFFF7FFFBFE07FFFFFFF33FFFFFFFE7100210EFFF7;
defparam prom_inst_29.INIT_RAM_2C = 256'h7FFFFFFD27FFFFFFFFBC0180037F9DCFFFFFE000106FFFFD7BD4FFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2D = 256'hFFFC004C60FFFFFEE7FFFFFFFFFFFFFFFFFFFFFFFFFD0C63FFFFFFFFFFFFDFE0;
defparam prom_inst_29.INIT_RAM_2E = 256'hFFFFFFFFFECE71FFFFFFFFFBFFFFF07FFFFFFC2FFFFFFFFFD31FFFCC1FFF7DFF;
defparam prom_inst_29.INIT_RAM_2F = 256'hFFFA5FFFFFFFFFDEFFFFFFFBCFFDFFFFFF81B0501FFFFFEFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_30 = 256'hF0000833FFFF5DFFFFFFFFFFFFFFFFFFFFFFFFFFE9B8FFFFFFFFFE7FEFE07FFF;
defparam prom_inst_29.INIT_RAM_31 = 256'hFFFFFFE4C63FFFFFFFFFFFE7F23FFFFFF8DFFFFFFFFFF7FFFFFFFF86EFFFFFFF;
defparam prom_inst_29.INIT_RAM_32 = 256'h3FFFFFFFFFFFFFFFFFFFFCDEBFFFFFFE0026307FFFF60E7FFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_33 = 256'hD8080FFFFF92DFFFFFFFFFFFFFFFFFFFFFFFFA231FFFFFFFFFF9E7F03FFFFFF4;
defparam prom_inst_29.INIT_RAM_34 = 256'hFFFBFB8FFFFFFFFFFF87FD1FFFFFF9BFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFC0;
defparam prom_inst_29.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFF97AF7FFFFF8000419FFFFBF77FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_36 = 256'h183FFFF9DFFFFFFFFFFFFFFFFFFFFFFFF900E7FFFFFFFFFFFFFC1FFFFFF07FFF;
defparam prom_inst_29.INIT_RAM_37 = 256'hC033FFFFFFFFFFFFFE0FFFFFF97FFFFFFFFFFFFFFFFFFFFFFF43DFFFFFFF0012;
defparam prom_inst_29.INIT_RAM_38 = 256'hFFFFEFFFFFFFFFFFF0FFFFFFFFF0680507FFFFFFFFFFFFFFFFFFFFFFFFFFFFFD;
defparam prom_inst_29.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9738FFFFFFFFFFFFFF87FFFFF97FFFFFFF;
defparam prom_inst_29.INIT_RAM_3A = 256'h7FFFFFFFFFFFFFC3FFFFF17FFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFC000004;
defparam prom_inst_29.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFE3BFFFFFFFC019041FFFFFFFFFFFFFFFFFFFFFFFFFFFFF99DC;
defparam prom_inst_29.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE8A33FFFFFFFFFFFFFC1FFFFF9FFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_3D = 256'hFFFFFFFFFFF4FFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF8340083FF;
defparam prom_inst_29.INIT_RAM_3E = 256'hFFFFFFFFFFFF3FFFFFFFFF0404827FFFF7FFFFFFFFFFFFFFFFFFFFFFEA618FFF;
defparam prom_inst_29.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFF49947FFFFFFFFFFFFF87FFFF97FFFFFFFFFFFFFDF;

pROM prom_inst_30 (
    .DO({prom_inst_30_dout_w[30:0],prom_inst_30_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_30.READ_MODE = 1'b1;
defparam prom_inst_30.BIT_WIDTH = 1;
defparam prom_inst_30.RESET_MODE = "SYNC";
defparam prom_inst_30.INIT_RAM_00 = 256'hFFFFFFFC3FFFFC3FFFFFFFFFFFFFF37FFFFFFFFFFFEFFFFFFFFFE00C2307FFFF;
defparam prom_inst_30.INIT_RAM_01 = 256'hFFFFFFFFFC3BFFFFFFFC0A8000FFFFFFFFFFFFFFFFFFFFFFFFFFFC7E33FFFFFF;
defparam prom_inst_30.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFE0618FFFFFFFFFFFFFE1FFFFE7FFFFFFFFFFFFFFDFFFF;
defparam prom_inst_30.INIT_RAM_03 = 256'hFFFF8FFFFF2FFFFFFFFFFFFFFF3FFFFFFFFFFFFF9FFFFFFFFF8202419FFFFFFF;
defparam prom_inst_30.INIT_RAM_04 = 256'hFFFFFFE3FFFFFFFFF0021127FFFFFFFFFFFFFFFFFFFFFFFFFF321C7FFFFFFFFF;
defparam prom_inst_30.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFC36B3FFFFFFFFFFFFF93FFFF97FFFFFFFFFFFFFF85FFFFFF;
defparam prom_inst_30.INIT_RAM_06 = 256'hE9FFFFEBFFFFFFFFFFFFFFE1DFFFFFFFFFFFF82FFFFFFFFE054040FFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_07 = 256'hFFFF0EFFFFFFFFC180205FFFFFFFFFFFFFFFFFFFFFFFFFDD718FFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_08 = 256'hFFFFFFFFFFFFE1F0C7FFFFFFFFFFFFF0FFFFE1FFFFFFFFFFFFFFFE7FFFFFFFFF;
defparam prom_inst_30.INIT_RAM_09 = 256'hFFF8FFFFFFFFFFFFFFFF9FFFFFFFFFFFFFE3DFFFFFFFFC010011FFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_0A = 256'hF87FFFFFFFFF8000283FFFFFFFFFFFFFFFFFFFFFFFF518E3FFFFFFFFFFFFF87F;
defparam prom_inst_30.INIT_RAM_0B = 256'hFFFFFFFFFE3918FFFFFFFFFFFFFE3FFFFC3FFFFFFFFFFFFFFFE5FFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_0C = 256'h1FFFFFFFFFFFFFFFF807FFFFFFFFFFFF0FFFFFFFFFF0C05007FFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_0D = 256'hFFFFFFFFFE00020CFFFFFFFFFFFFFFFFFFFFFFFE8B8C7FFFFFFFFFFFFE4FFFFF;
defparam prom_inst_30.INIT_RAM_0E = 256'hFFFFFF8F863FFFFFFFFFFFFF87FFFFAFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFC3;
defparam prom_inst_30.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFE3BFFFFFFFFFFFFBFFFFFFFFFFC009041FFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_10 = 256'hFFFFFFF8441903FFFFFFFFFFFFFFFFFFFFFFB0C58FFFFFFFFFFFFFC3FFFF87FF;
defparam prom_inst_30.INIT_RAM_11 = 256'hFF03D8C7FFFFFFFFFFFFE1FFFFE9FFFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_12 = 256'hFFFFFFFFFFFE06FFFFFFFFFFFFBFFFFFFFFFFF0001043FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_13 = 256'hFFFFE0144407FFFFFFFFFFFFFFFFFFFC0F1063FFFFFFFFFFFFF87FFFF8FFFFFF;
defparam prom_inst_30.INIT_RAM_14 = 256'h5E58FFFFFFFFFFFFFC3FFFFC3FFFFFFFFFFFFFFFFFC1DFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_15 = 256'hFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFC0B0440FFFFFFFFFFFFFFFFFC4084;
defparam prom_inst_30.INIT_RAM_16 = 256'hFFE40001BFFFFFFFFFFFFFFFF87002C6AC3FFFFFFFFFFFFE5FFFFC1FFFFFFFFF;
defparam prom_inst_30.INIT_RAM_17 = 256'h0FFFFFFFFFFFFF87FFFFCFFFFFFFFFFFFFFFFFFF00BFFFFFFFFFFEFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_18 = 256'hFFFFFFE027FFFFFFFFFE3FFFFFFFFFFFF0025183FFFFFFFFFFFFFFFDF8538EC6;
defparam prom_inst_30.INIT_RAM_19 = 256'h8C40007FFFFFFFFFFFFFFCFD381A4587FFFFFFFFFFFFE3FFFF87FFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_1A = 256'hFFFFFFFFFFE5FFFFC9FFFFFFFFFFFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_30.INIT_RAM_1B = 256'hFFFFC07FFFFFFFFFFFFFFFFFFFFFFFD301204FFFFFFFFFFFFFFE87F82992E1FF;
defparam prom_inst_30.INIT_RAM_1C = 256'h2811FFFFFFFFFFFFFF1F8C3129303FFFFFFFFFFFF87FFFF4FFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_1D = 256'hFFFFFFFCBFFFFC7FFFFFFFFFFFFFFFFFFFF009FFFFFFFFF3FFFFFFFFFFFFFE01;
defparam prom_inst_30.INIT_RAM_1E = 256'hFE237FFFFFFFFFFFFFFFFFFFFFFFC0A0083FFFFFFFFFFFFFBFC413C8E607FFFF;
defparam prom_inst_30.INIT_RAM_1F = 256'h07FFFFFFFFFFFFEFF00F337F41FFFFFFFFFFFF0FFFFE1FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_20 = 256'hFFFF97FFFF0FFFFFFFFFFFFFFFFFFFFFE001FFFFFF01FFFFFFFFFFFFFFE84054;
defparam prom_inst_30.INIT_RAM_21 = 256'h0021FFFE8CDFFFFFFFFFFFFFFD001204FFFFFFFFFFFFFFDC0F11DFE83FFFFFFF;
defparam prom_inst_30.INIT_RAM_22 = 256'hFFFFFFFFFFFDEE1F7FCFF907FFFFFFFFFFE1FFFFD3FFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_30.INIT_RAM_23 = 256'hF2FFFFF1FFFFFFFFFFFFFFFFFFFFFF840021C60187FFFFFFFFFFFFFFE00A041F;
defparam prom_inst_30.INIT_RAM_24 = 256'h00001803FFFFFFFFFFFFFFF47A12A3FFFFFFFFFFFF7B9F13E3FF61FFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_25 = 256'hFFFFFFFF978F01D8FFCC3FFFFFFFFFFEBFFFF27FFFFFFFFFFFFFFFFFFFFFF800;
defparam prom_inst_30.INIT_RAM_26 = 256'hFFFE3FFFFFFFFFFFFFFFFFFFFFFF8000218207FFFFFFFFFFFFFFFE8009043FFF;
defparam prom_inst_30.INIT_RAM_27 = 256'h0007FFFFFFFFFFFFFFFFD014068FFFFFFFFFFFC587C04F7FFB0FFFFFFFFFFF1F;
defparam prom_inst_30.INIT_RAM_28 = 256'hFFFFF1C1E077E79CA3FFFFFFFFFF97FFFF5FFFFFFFFFFFFFFFFFFFF1DFF02000;
defparam prom_inst_30.INIT_RAM_29 = 256'h87FFFFFFFFFFFFFFFFFFFBFB7FF020001FFFFFFFFFFFFFFFFFFE140161FFFFFF;
defparam prom_inst_30.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFF4204803FFFFFFFFFFC10E015F3FF38FFFFFFFFFFE3FFFF;
defparam prom_inst_30.INIT_RAM_2B = 256'hFF003C0ABCFFC63FFFFFFFFFF0FFFFE1FFFFFFFFFFFFFFFFFFF9FFCFFFF0008F;
defparam prom_inst_30.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFF4BFFCBFFFFFFFFFFFFFFFFFFFFFFFFFC800100FFFFFFFFF;
defparam prom_inst_30.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFD005401FFFFFFFFFF180F8057FFF48FFFFFFFFFFCFFFFF0FF;
defparam prom_inst_30.INIT_RAM_2E = 256'h8381F7BFF823FFFFFFFFFF1FFFFE3FFFFFFFFFFFFFFFFFE7DFFFEBFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_2F = 256'hFFFFFFFFFFFFE33FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFA75000FFFFFFFFFF81;
defparam prom_inst_30.INIT_RAM_30 = 256'hFFFFFFFFFFFFFC40003FFFFFFFFFEB60FEBBFFFEB9FFFFFFFFFF87FFFF0FFFFF;
defparam prom_inst_30.INIT_RAM_31 = 256'hD6FFFF447FFFFFFFFFE7FFFF83FFFFFFFFFFFFFFFFE1DFFFFFEBFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_32 = 256'hFFFFFFFFE0EF7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFD800007FFFFFFFFDEC01E;
defparam prom_inst_30.INIT_RAM_33 = 256'hFFFFFFFFFFF00003FFFFFFFF999807E1FFFF831FFFFFFFFFFCFFFFE1FFFFFFFF;
defparam prom_inst_30.INIT_RAM_34 = 256'hFF828FFFFFFFFFFE3FFFFC7FFFFFFFFFFFFFFFF0D7FBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_35 = 256'hFFFFF06BFFBFFFCF7FFFFFFFFFFFFFFFFFFFFFFFF30001FFFFFFFF980E307FFB;
defparam prom_inst_30.INIT_RAM_36 = 256'hFFFFFFFE80007FFFFFFF98057822F2FFC143FFFFFFFFFFCFFFFF1FFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_37 = 256'hB1FFFFFFFFFFCFFFFFA7FFFFFFFFFFFFFFF804FFFBFFFDFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_38 = 256'hFE0C7FFF3FFF1DFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFC87AF6DEEFFFC4;
defparam prom_inst_30.INIT_RAM_39 = 256'hFFFFFE805FFFFFFFC817BFF75CFFE258FFFFFFFFFFF3FFFFE1FFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3A = 256'hFFFFFFFFFC7FFFFAFFFFFFFFFFFFFFFE023FFFF3FFF3EFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3B = 256'h9FFFF13FFE5EFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFFFC100F1DFFF7FF00C7F;
defparam prom_inst_30.INIT_RAM_3C = 256'hFFFFFFFFFFFFF0F0D8DFEAFFF9063FFFFFFFFFFE1FFFFC3FFFFFFFFFFFFFFF03;
defparam prom_inst_30.INIT_RAM_3D = 256'hFFFFFF97FFFF07FFFFFFFFFFFFFF81EFFFF013FFD9FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3E = 256'hFC011FF89FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0300E1EFD5FFE971FFFFF;
defparam prom_inst_30.INIT_RAM_3F = 256'hFFFFFFFFF80C4381FABFFE4B8FFFFFFFFFFFF7FFFFE3FFFFFFFFFFFFFF8073FF;

pROM prom_inst_31 (
    .DO({prom_inst_31_dout_w[30:0],prom_inst_31_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_31.READ_MODE = 1'b1;
defparam prom_inst_31.BIT_WIDTH = 1;
defparam prom_inst_31.RESET_MODE = "SYNC";
defparam prom_inst_31.INIT_RAM_00 = 256'hFFFFFFF6CE120000000000000000400000009860000000000000000000000003;
defparam prom_inst_31.INIT_RAM_01 = 256'h40000000000000000000000000000040000000000000000000000000047FFFFF;
defparam prom_inst_31.INIT_RAM_02 = 256'h000000000000000000000009FFFFFFFFFFFFFFBFC08100008980020078240000;
defparam prom_inst_31.INIT_RAM_03 = 256'hFFFFDEA680000000000003004580000023924000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_04 = 256'h182228000000000000000000000000000000000000000000000001EFFFFF97FF;
defparam prom_inst_31.INIT_RAM_05 = 256'h000000000000000000013FFFFF9F7FFFFFFFFEC682000600000037E609E27FF8;
defparam prom_inst_31.INIT_RAM_06 = 256'hFFFFE7B10801860000CFFDEFFF9FFE6665890000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_07 = 256'h1F0300000000000000000000000000000000000000000000012FFFFFCFF7FFFF;
defparam prom_inst_31.INIT_RAM_08 = 256'h0000000000000041BFFFFFCFFF1FFFFFFFFDE486200000B3FDF7EFFEF7FCD4BC;
defparam prom_inst_31.INIT_RAM_09 = 256'hFEFF9C804BE179FFFFFFBFBFF499B5D2FD300000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_0A = 256'h400000000000000000000000000000000000000000004DF7FFFFAFFFF3FFFFFF;
defparam prom_inst_31.INIT_RAM_0B = 256'h000000000010BDFFFFE7FFFF3FFFFFFFA7E70017F85F7FFFF7DFAFFD3795779F;
defparam prom_inst_31.INIT_RAM_0C = 256'hFE007969FFCFF7DFFFFFFFEFB63FFD8000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000008BFFFFF3FFFF00FFFFFFFF;
defparam prom_inst_31.INIT_RAM_0E = 256'h0000000004FFFFF83FFF839FFFFEF7FF801FDF7FF3FEFFFFFFFFFFE57FFFC800;
defparam prom_inst_31.INIT_RAM_0F = 256'h01F97FFFFFFDFFFFFFFFE7B1F7E0000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_10 = 256'h000000000000000000000000000000000000010CBFFFF303FF83F9FFFFFFDBE0;
defparam prom_inst_31.INIT_RAM_11 = 256'h000002FF7FFBF03F81FF8FFFEFFAC60879BBF3FFFFFFFFDFFFFC7510F2030000;
defparam prom_inst_31.INIT_RAM_12 = 256'h6EFCFFFFFFFFFFFFFF9DD23E0000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_13 = 256'h000000000000000000000000000000000044BFBFF3FF03C1FFF95FBEFF30041E;
defparam prom_inst_31.INIT_RAM_14 = 256'h005BFFF1FFF001FFFF9FF8060180247C8FFFFFFFFFFFEF7FFF62E38C00000000;
defparam prom_inst_31.INIT_RAM_15 = 256'hEFFFF3FFFFF7FFFFFE7BB0A00000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_16 = 256'h0000000000000000000000000000000001FFF1FFFF08FFFFE2C008200002069D;
defparam prom_inst_31.INIT_RAM_17 = 256'h7FFCFFFFE03FFFF0400000000110077FFF0FFFFFFFFFFFFFBD13A01000101000;
defparam prom_inst_31.INIT_RAM_18 = 256'hFDBFFE7EFFFFFFFF070002000010000000000000000000000000000000000010;
defparam prom_inst_31.INIT_RAM_19 = 256'h00000000000000000000000000000497FA7FFFE003FFF87C000000100085FFFF;
defparam prom_inst_31.INIT_RAM_1A = 256'h0FFFF0303FF83FC000100000193FFFFFFFFF97BFFFFF9FDDCC00004000400000;
defparam prom_inst_31.INIT_RAM_1B = 256'hFFFF7FFFFFFFC2C0250000000000000000000000000000000000000000013BFF;
defparam prom_inst_31.INIT_RAM_1C = 256'h000000000000000000000000040ED8407FF03F03F83FFC02000000019FFFFFFF;
defparam prom_inst_31.INIT_RAM_1D = 256'hF83FF03C1FFFC4000000001FFFFFFFFEFEFEFFFFFFF4F1003000000080000000;
defparam prom_inst_31.INIT_RAM_1E = 256'h3F5FFFFFFD3C00202010002000000000000000000000000000000000149F7C07;
defparam prom_inst_31.INIT_RAM_1F = 256'h0000000000000000000000040E7FC0781FFF001FFFFC0000000007FFFFFF00FE;
defparam prom_inst_31.INIT_RAM_20 = 256'hFFF00FFFFE0000000089E7FFF400CEBFFFAAFFDFDF0050000800000000000000;
defparam prom_inst_31.INIT_RAM_21 = 256'hFEFFFFB06820000000008000000000000000000000000000000010033FFC001F;
defparam prom_inst_31.INIT_RAM_22 = 256'h00000000000000000000403FFFC00FFFFE00FFFF000000000B7FFFFA03FC7DFF;
defparam prom_inst_31.INIT_RAM_23 = 256'h000FFF0000000009BFFFFE0FF883FFFFDAFEFCF8040004000000000000000000;
defparam prom_inst_31.INIT_RAM_24 = 256'hBFFE9020240000000400000000000000000000000000000000041FFFFC07FFFF;
defparam prom_inst_31.INIT_RAM_25 = 256'h00000000000000000C1FFFFE10FFFF8381FF8000000000BFFFFC1FDFDA7FFFFF;
defparam prom_inst_31.INIT_RAM_26 = 256'h1F8200000001B7FFFC1FDA1B1FFFFFEFFD960806040200100008000000000000;
defparam prom_inst_31.INIT_RAM_27 = 256'hFFF002000884C0180000000000000000000000000000000327FFFE000FFF83F8;
defparam prom_inst_31.INIT_RAM_28 = 256'h00000000000000107FFF0780FF81FF81C0000000000FFFDF8FFE83E1FFFFFBFF;
defparam prom_inst_31.INIT_RAM_29 = 256'h00000000037FFFC3F867F11FFFFFFFFFF1200043032680000000000000000000;
defparam prom_inst_31.INIT_RAM_2A = 256'h780000C0CC20000200000000000000000000000000000007FF03FC0FC0FFF801;
defparam prom_inst_31.INIT_RAM_2B = 256'h000000000000B07F81FFC0C0FFFF800000000002DFFFE0F80DC001FFFFFFFFFC;
defparam prom_inst_31.INIT_RAM_2C = 256'h0000005FFFF81E0F80006FFFFFFFFFE110018008460004000000000000000000;
defparam prom_inst_31.INIT_RAM_2D = 256'h0C0000401120000000000000000000000000000000010781FFFC007FFFF04000;
defparam prom_inst_31.INIT_RAM_2E = 256'h00000000021000FFFFC07FFFF8000000000029FFBC03FF000003FFFFFFFFFFC3;
defparam prom_inst_31.INIT_RAM_2F = 256'h0019FDFF007B000000FFFFFFFFFFF3C1802422040E0000000000000000000000;
defparam prom_inst_31.INIT_RAM_30 = 256'h48010011000200000000000000000000000000000100FFFFF18FFFFC30000000;
defparam prom_inst_31.INIT_RAM_31 = 256'h00000010107FFFF8007FFC250080000002BFFFC00E8000080FFFFFFFFFFF40C0;
defparam prom_inst_31.INIT_RAM_32 = 256'h2FDFC00100001B02FFFFA77FFFE0300019410420000000000000000000000000;
defparam prom_inst_31.INIT_RAM_33 = 256'h61018000080000000000000000000000000000020FFFF8100FFE114040000000;
defparam prom_inst_31.INIT_RAM_34 = 256'h00008000FFFC1FC07E00504000000007FFFE80200003E07FFFE215FEFFB20004;
defparam prom_inst_31.INIT_RAM_35 = 256'hFFE80400E3FC07FFF7FFEF7F3C110A6803000100040000000000000000000000;
defparam prom_inst_31.INIT_RAM_36 = 256'h9E9802000000000000000000000000000020060FFC0FFC07080424000000003F;
defparam prom_inst_31.INIT_RAM_37 = 256'h000420FE0FFFC0000100000000000FFFB80000E62781FFFA7FF9DBCC07401C01;
defparam prom_inst_31.INIT_RAM_38 = 256'h0020EF8FD85FFFD9FDFFD9230204080320800400000000000000000000000000;
defparam prom_inst_31.INIT_RAM_39 = 256'h0001000000000000000000000000000081220E07FFFC0400100000000223D7B0;
defparam prom_inst_31.INIT_RAM_3A = 256'h082007FFFF8000410000000000A28C00041F9C9F07FFFFFFDFFE5C8000B00050;
defparam prom_inst_31.INIT_RAM_3B = 256'hF39F3FE0FFFFFFFFDFC800101880581894C00000000000000000000000000008;
defparam prom_inst_31.INIT_RAM_3C = 256'h0200000000000000000000000000098A0203FFFFC20010000000000000220000;
defparam prom_inst_31.INIT_RAM_3D = 256'h00FFFFE18004000000000000000000077E733C0FFFFFFFFFA7330001E61891E4;
defparam prom_inst_31.INIT_RAM_3E = 256'h7C7F83FFFFFFFFD9CCC0006186261C0080000000000000000000000000039840;
defparam prom_inst_31.INIT_RAM_3F = 256'h000000000000000000000000000990000FFFE10003200000000000000000006F;

pROM prom_inst_32 (
    .DO({prom_inst_32_dout_w[30:0],prom_inst_32_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_32.READ_MODE = 1'b1;
defparam prom_inst_32.BIT_WIDTH = 1;
defparam prom_inst_32.RESET_MODE = "SYNC";
defparam prom_inst_32.INIT_RAM_00 = 256'hFFF08001000000000000000200000DFCECB03FFFFF7FF4BF010A0781BBDCCEB0;
defparam prom_inst_32.INIT_RAM_01 = 256'hFE0FFFFFFFFFC8010040181C06C2880000000000000000000000000014800100;
defparam prom_inst_32.INIT_RAM_02 = 256'h00000000000000000000000011804A0FF802011400000000000010000001BDF1;
defparam prom_inst_32.INIT_RAM_03 = 256'h40D0900000000000000004000037F3F2E0FFFFFFFFFB006014860E9841009000;
defparam prom_inst_32.INIT_RAM_04 = 256'h1FFFFFFF7B714200000FC78820200000000000000000000000000001300020F8;
defparam prom_inst_32.INIT_RAM_05 = 256'h00000000000000000000202100020C00140000A0000000026000040007FBE3FC;
defparam prom_inst_32.INIT_RAM_06 = 256'hC00050000000010000000800FFE7ED81FFFFFFFDDC9088608478C00600000000;
defparam prom_inst_32.INIT_RAM_07 = 256'hFFFFFFFEA0002101BF7E8100000000000000000000000000000000A290202004;
defparam prom_inst_32.INIT_RAM_08 = 256'h0000000000000000000102000210010400300000000000000000000FEF8BF01F;
defparam prom_inst_32.INIT_RAM_09 = 256'h28000000004007F8000001FF93F603FFFFFFFFC0020000069800000000000000;
defparam prom_inst_32.INIT_RAM_0A = 256'hFFF3C000000019E7800000000000000000000000000000002049200004000000;
defparam prom_inst_32.INIT_RAM_0B = 256'h0000000000000002021320090002001400000000001F018000003FE727C07FFF;
defparam prom_inst_32.INIT_RAM_0C = 256'h000000000C000E000007FFCFF80FDFFFFFD20000071FEE068721000000000000;
defparam prom_inst_32.INIT_RAM_0D = 256'hEC00206180E512E0008000000000000000000200000000220108020004000000;
defparam prom_inst_32.INIT_RAM_0E = 256'h210081000000A29003000000000000000000000C0000700000FFDECF00BFFEFF;
defparam prom_inst_32.INIT_RAM_0F = 256'h00020400000380001FDF1FE00FFFFFFF60080020608758100000000000000000;
defparam prom_inst_32.INIT_RAM_10 = 256'h200002185F072200000000000000000000204048000200020000048804800000;
defparam prom_inst_32.INIT_RAM_11 = 256'h001000000420000200825A00202000000003000000300003FF3F2C0004FFFC20;
defparam prom_inst_32.INIT_RAM_12 = 256'h008000000300007F7E7FC001BDFF000B00010006F0C8A0000000000000000404;
defparam prom_inst_32.INIT_RAM_13 = 256'h00000C7B80820000000000000001010004102000002004210246822810000000;
defparam prom_inst_32.INIT_RAM_14 = 256'h040800204805020120A14A08000000004000000040000FFEDED8002FDC302101;
defparam prom_inst_32.INIT_RAM_15 = 256'h000000080201FFB89F1F81330C08000000196EE7010000000000000030404042;
defparam prom_inst_32.INIT_RAM_16 = 256'h06CDB7E000000000000000208810048102000808410431002022800000000810;
defparam prom_inst_32.INIT_RAM_17 = 256'h000002044040100080A400000000080000000180003FBF3F00000CC10001200C;
defparam prom_inst_32.INIT_RAM_18 = 256'h0000302007FE7F0000000000CA06030110431000000000000000000000012021;
defparam prom_inst_32.INIT_RAM_19 = 256'h8F84000000000000000004002044190000005442040000103A00000001020000;
defparam prom_inst_32.INIT_RAM_1A = 256'h041444804000C808000000004080000000040000FE7F000000400304040007A6;
defparam prom_inst_32.INIT_RAM_1B = 256'h0180001FFF807000040001080021819FC01000000000000000004000100C0000;
defparam prom_inst_32.INIT_RAM_1C = 256'h0420000000000000000400000000000040000000001403000000001000000000;
defparam prom_inst_32.INIT_RAM_1D = 256'hA0000240110080000000060000000000200003FF80600000004120081E04457D;
defparam prom_inst_32.INIT_RAM_1E = 256'h00007E0040000008004403662168AFCF0800000000000001C038000000000004;
defparam prom_inst_32.INIT_RAM_1F = 256'h0000000000000000000000020000006808808000404000000000810000000008;
defparam prom_inst_32.INIT_RAM_20 = 256'h00000950200000000020400000000200000E0000000001000010040060B0E788;
defparam prom_inst_32.INIT_RAM_21 = 256'h0190000000002000412007782674000000000000000000800000008000000701;
defparam prom_inst_32.INIT_RAM_22 = 256'h0000000000000000000000000000400080041800000000000800000000008000;
defparam prom_inst_32.INIT_RAM_23 = 256'h0006100000000003010000000020400030000000000000024001DE19F7000000;
defparam prom_inst_32.INIT_RAM_24 = 256'h0000000000000018007A02170FC0000000000000000100000000000000040891;
defparam prom_inst_32.INIT_RAM_25 = 256'h0000000000000000038000000082494A41880000000000600000000010100006;
defparam prom_inst_32.INIT_RAM_26 = 256'h240000000000080000000000000001C000000000200000000001F1ECB2000000;
defparam prom_inst_32.INIT_RAM_27 = 256'h000000000002000860185E020000000000000000020000002000000008909020;
defparam prom_inst_32.INIT_RAM_28 = 256'h0000000000000004000000008400000000000000000200000000040400007000;
defparam prom_inst_32.INIT_RAM_29 = 256'h000000000040000000000200000800000000010000000A1667F7D00000000000;
defparam prom_inst_32.INIT_RAM_2A = 256'h00000000005EE399CCF8A0000000000000000000000000800000000C00000000;
defparam prom_inst_32.INIT_RAM_2B = 256'h00000000000000000000000010010000000000001C0800000000000006000000;
defparam prom_inst_32.INIT_RAM_2C = 256'h0000000302000000804000010000000000000000019700BB972E000000000000;
defparam prom_inst_32.INIT_RAM_2D = 256'h0000000007094ABE118000000000000000000000000400000000080400800000;
defparam prom_inst_32.INIT_RAM_2E = 256'h0008000000800000000001004000000000000040400000006000006000000000;
defparam prom_inst_32.INIT_RAM_2F = 256'h0000180000000010000018000000000000000041C49487860000000000000000;
defparam prom_inst_32.INIT_RAM_30 = 256'h000600058A7D7E08000000000000000000000000200000000010084000000000;
defparam prom_inst_32.INIT_RAM_31 = 256'h0000000400000000010820000000000000030000000008000007000000000000;
defparam prom_inst_32.INIT_RAM_32 = 256'h00404430000C000001C000000000000000008281F829C8000000000000000000;
defparam prom_inst_32.INIT_RAM_33 = 256'h0041E0D201BA0000000000000000000000000100000000001210000000000000;
defparam prom_inst_32.INIT_RAM_34 = 256'h00004000000000019800000000000000100000001C0000003800000000000000;
defparam prom_inst_32.INIT_RAM_35 = 256'h000000180000000700000000010000000780EE62680000000000000000000800;
defparam prom_inst_32.INIT_RAM_36 = 256'h01BC711640000000000000000000000000300000000000000000000000000002;
defparam prom_inst_32.INIT_RAM_37 = 256'h0800000000000000000000000000007400083800000000E00100000100000060;
defparam prom_inst_32.INIT_RAM_38 = 256'h0230000000003C0000000080000000E04296F400000000000000000000400000;
defparam prom_inst_32.INIT_RAM_39 = 256'hF3BDC0C000000000000000000000000600000000000000000000000000000780;
defparam prom_inst_32.INIT_RAM_3A = 256'h000000000000000000000000000030C1F0000000000780000000000000000018;
defparam prom_inst_32.INIT_RAM_3B = 256'h0000040000F00000000000000000003EEF3000000000000000000002000003C0;
defparam prom_inst_32.INIT_RAM_3C = 256'hF500000000000000000000C00001F0000000000000000000000000000007FFD0;
defparam prom_inst_32.INIT_RAM_3D = 256'h00000000000000000000000000001000000000000E00000000000000001E71AF;
defparam prom_inst_32.INIT_RAM_3E = 256'h00740001C0000001000000440F41BEFF280000000000000000000000037E0000;
defparam prom_inst_32.INIT_RAM_3F = 256'h000000000000000000010017EF80000000000000000000000000000000000000;

pROM prom_inst_33 (
    .DO({prom_inst_33_dout_w[30:0],prom_inst_33_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_33.READ_MODE = 1'b1;
defparam prom_inst_33.BIT_WIDTH = 1;
defparam prom_inst_33.RESET_MODE = "SYNC";
defparam prom_inst_33.INIT_RAM_00 = 256'h0000000000000000000000000000000045000038000001FE0000100241D7BFE0;
defparam prom_inst_33.INIT_RAM_01 = 256'h000007800001FF80000041839813D000000000000000000000087FFDC0000000;
defparam prom_inst_33.INIT_RAM_02 = 256'h000000000000000000BFFFF00000000000000000000000000000000000000218;
defparam prom_inst_33.INIT_RAM_03 = 256'h0000000000000000000000000000470000007E0003FFF000010A031A3C799000;
defparam prom_inst_33.INIT_RAM_04 = 256'h0007FC41FFF6000183045FDB21200000000000000000000015F8F80000000000;
defparam prom_inst_33.INIT_RAM_05 = 256'h0000000000000000F07C00000000000000000000000000000000000000003100;
defparam prom_inst_33.INIT_RAM_06 = 256'h00000000000000000000000000440000000F987FE7C0000000183B841E000000;
defparam prom_inst_33.INIT_RAM_07 = 256'h00327FC7F80006000E0F000B8000000000000000000000263F00000000000000;
defparam prom_inst_33.INIT_RAM_08 = 256'h0000000000000CFF000000000000000000000000000000000000000001000000;
defparam prom_inst_33.INIT_RAM_09 = 256'h00000000000000000000000800000000023F91FB00006200319CFD0000000000;
defparam prom_inst_33.INIT_RAM_0A = 256'h7FB7F3E0008000E077B7800000000000000000000001FF000000000000000000;
defparam prom_inst_33.INIT_RAM_0B = 256'h0000000000180000000000000000000000000000000000000000004600000000;
defparam prom_inst_33.INIT_RAM_0C = 256'h0000000000000000003010000000000DFFE3FC0000002005EBF3000000000000;
defparam prom_inst_33.INIT_RAM_0D = 256'hC8EF80064800041F8A0000000000000000000000000000000000000000000000;
defparam prom_inst_33.INIT_RAM_0E = 256'h00000000000000000000000000000000000000000000000300000000000001BF;
defparam prom_inst_33.INIT_RAM_0F = 256'h000000000000000000040000000037D3F9F01214238107D98000000000000000;
defparam prom_inst_33.INIT_RAM_10 = 256'hF600010E0000D7A0000000000000000000000000000000000000000000000000;
defparam prom_inst_33.INIT_RAM_11 = 256'h000000000180000000000000000000000000000000070080000400000003FFF1;
defparam prom_inst_33.INIT_RAM_12 = 256'h000000001FFC000000000000007FE477C004000058D400000000000000000000;
defparam prom_inst_33.INIT_RAM_13 = 256'h0110001619F80000000000000000000000000000040000000000000000000000;
defparam prom_inst_33.INIT_RAM_14 = 256'h000000180000000000000000000000000000007E00000000000000000FC9FCF8;
defparam prom_inst_33.INIT_RAM_15 = 256'h0007F8000000000000000001FFF1FB00610099610C0000000000000000000000;
defparam prom_inst_33.INIT_RAM_16 = 256'h001899C360000000000000000000000000000E20000000000000000000000000;
defparam prom_inst_33.INIT_RAM_17 = 256'h000B1800000000000000000000000000FFC00000000000000000003FE27BE006;
defparam prom_inst_33.INIT_RAM_18 = 256'h0000000000000000000007E5F67C0400000451E4000000000000000000000000;
defparam prom_inst_33.INIT_RAM_19 = 256'h0109280000000000000000000000000001842000000040020000000000007FFC;
defparam prom_inst_33.INIT_RAM_1A = 256'hE508000000000010000000000FFC000000000000000000000000FFF8FD801000;
defparam prom_inst_33.INIT_RAM_1B = 256'h0000000000000000001FF139F004000A26590000000000000000000000000002;
defparam prom_inst_33.INIT_RAM_1C = 256'h0120000000000000000000000000015382000000100000000000003F00000000;
defparam prom_inst_33.INIT_RAM_1D = 256'h80000000000010000000FC0000000000000000000000000003F6FB7E01000000;
defparam prom_inst_33.INIT_RAM_1E = 256'h00000000000000007FFC7EC00000032682000000000000000000000000009943;
defparam prom_inst_33.INIT_RAM_1F = 256'h800000000000000000000000002CA0C0000002000000000001F0000000000000;
defparam prom_inst_33.INIT_RAM_20 = 256'h0000800000800003E0000000000000000001C0000000000FF99CF800000149B4;
defparam prom_inst_33.INIT_RAM_21 = 256'h38000000000001FB7DBF0000002000000000000000000000000000000B727000;
defparam prom_inst_33.INIT_RAM_22 = 256'h0000000000000000000000001938000000200000200007C00000000000FF0000;
defparam prom_inst_33.INIT_RAM_23 = 256'h08000000000F8000000000400000000003C0000000003FFE3E60000004843000;
defparam prom_inst_33.INIT_RAM_24 = 256'h000000000007FCCE7C000004013000000000000000000000000001000C000000;
defparam prom_inst_33.INIT_RAM_25 = 256'h00000000000000000000B00600000002000004000F00000000080F000000003C;
defparam prom_inst_33.INIT_RAM_26 = 256'h0000001E0000000001C00000000000000000000000F9BEDF8000008040000000;
defparam prom_inst_33.INIT_RAM_27 = 256'h000000001FFF1F300000086F0000000000000000000000000001870000000000;
defparam prom_inst_33.INIT_RAM_28 = 256'h0000000000000000000700000000100001001C00000000060000000000000000;
defparam prom_inst_33.INIT_RAM_29 = 256'h801C000000001800000000000000001000200003FE673E000000C44000000000;
defparam prom_inst_33.INIT_RAM_2A = 256'h0000007CDE6FC000021180000000000000000000000000080380000000040000;
defparam prom_inst_33.INIT_RAM_2B = 256'h0000000000000401C0000000008000401C000000011000000000000000000008;
defparam prom_inst_33.INIT_RAM_2C = 256'h0000000020000000000000000000023000000FFF8F980002842B000000000000;
defparam prom_inst_33.INIT_RAM_2D = 256'h0001FF339F000001180000000000000000000000000000E0000000002000201C;
defparam prom_inst_33.INIT_RAM_2E = 256'h00000000000030000000000400101C0000000260000000000000000000008200;
defparam prom_inst_33.INIT_RAM_2F = 256'h00004000000000000000000000020000003E4FA7E00000100000000000000000;
defparam prom_inst_33.INIT_RAM_30 = 256'h07FFC7CC0000A2000000000000000000000000000418000000000080100C0000;
defparam prom_inst_33.INIT_RAM_31 = 256'h000000000E000000000020100E00000004400000000000000000000000000000;
defparam prom_inst_33.INIT_RAM_32 = 256'h80000000000000000000000040000000FF99CF800009F1800000000000000000;
defparam prom_inst_33.INIT_RAM_33 = 256'h27F3F000006D2000000000000000000000001007000000000006100600000000;
defparam prom_inst_33.INIT_RAM_34 = 256'h000801800000000000F00700000008800000000000000000000000000000001F;
defparam prom_inst_33.INIT_RAM_35 = 256'h000000000000000000000008000003FFE3E60000408800000000000000000000;
defparam prom_inst_33.INIT_RAM_36 = 256'hE7C000062000000000000000000000000004E000000000000003000000090000;
defparam prom_inst_33.INIT_RAM_37 = 256'h0270000000000000018000000100000000000000000000000000000000007FCC;
defparam prom_inst_33.INIT_RAM_38 = 256'h000000000000000000000000000F93F8F8000000000000000000000000000000;
defparam prom_inst_33.INIT_RAM_39 = 256'h000000000000000000000000000000001800000000000000C000000100000000;
defparam prom_inst_33.INIT_RAM_3A = 256'h0000000000000060000009000000000000000000000000000000000001FFF1FB;
defparam prom_inst_33.INIT_RAM_3B = 256'h0000000000000000000000003FE67BE00000000000000000000000000000400C;
defparam prom_inst_33.INIT_RAM_3C = 256'h0000000000000000000000000024070000000000000010000009000000000000;
defparam prom_inst_33.INIT_RAM_3D = 256'h00000000000C00000100000000000000000000000000000000000007C9FE7C00;
defparam prom_inst_33.INIT_RAM_3E = 256'h0000000000000000000000FBF87D800008000000000000000000000000138000;
defparam prom_inst_33.INIT_RAM_3F = 256'h00000000000000000000000000C0000000000000060000000000000000000000;

pROM prom_inst_34 (
    .DO({prom_inst_34_dout_w[30:0],prom_inst_34_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_34.READ_MODE = 1'b1;
defparam prom_inst_34.BIT_WIDTH = 1;
defparam prom_inst_34.RESET_MODE = "SYNC";
defparam prom_inst_34.INIT_RAM_00 = 256'h00000003000002800000000000000000000000000000000000001FF39CF00000;
defparam prom_inst_34.INIT_RAM_01 = 256'h00000000000000000003F47F3E00000000000000000000000000000070000000;
defparam prom_inst_34.INIT_RAM_02 = 256'h0000000000000000000101380000000000000180000140000000000000000000;
defparam prom_inst_34.INIT_RAM_03 = 256'h0000C00000A0000000000000000000000000000000000000007DFC3E40000000;
defparam prom_inst_34.INIT_RAM_04 = 256'h00000000000000000FFDCEDC00000000000000000000000000808C0000000000;
defparam prom_inst_34.INIT_RAM_05 = 256'h0000000000000000408700000000000000300000500000000000000000000000;
defparam prom_inst_34.INIT_RAM_06 = 256'h180000280000000000000000000000000000000000000001FA3F9F8000000000;
defparam prom_inst_34.INIT_RAM_07 = 256'h000000000000003E7F1FB0000000000000000000000000000380000000000000;
defparam prom_inst_34.INIT_RAM_08 = 256'h0000000000000009C00000000000000C00000400000000000000000000000000;
defparam prom_inst_34.INIT_RAM_09 = 256'h0002000000000000000000000000000000000000000007FEE7EE000000000000;
defparam prom_inst_34.INIT_RAM_0A = 256'h000000000000FF9FC7C000000000000000000000000204600000000000000600;
defparam prom_inst_34.INIT_RAM_0B = 256'h0000000000023800000000000003000000000000000000000000000000000000;
defparam prom_inst_34.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000001F3F8FF800000000000000;
defparam prom_inst_34.INIT_RAM_0D = 256'h0000000003FFF1F3000000000000000000000001001C00000000000000C00000;
defparam prom_inst_34.INIT_RAM_0E = 256'h000000804E00000000000000600000A000000000000000000000000000000000;
defparam prom_inst_34.INIT_RAM_0F = 256'h00000000000000000000000000000000000000007FC6F3E00000000000000000;
defparam prom_inst_34.INIT_RAM_10 = 256'h0000000F9BE6FC00000000000000000000000023800000000000003000001000;
defparam prom_inst_34.INIT_RAM_11 = 256'h000001C000000000000008000000000000000000000000000000000000000000;
defparam prom_inst_34.INIT_RAM_12 = 256'h00000000000000000000000000000000000001FFF8F980000000000000000000;
defparam prom_inst_34.INIT_RAM_13 = 256'h00003FE339F000000000000000000000000CE000000000000006000000000000;
defparam prom_inst_34.INIT_RAM_14 = 256'h2038000000000000030000040000000000000000000000000000000000000000;
defparam prom_inst_34.INIT_RAM_15 = 256'h000000000000000000000000000000000007E4FB3E000000000000000001FF80;
defparam prom_inst_34.INIT_RAM_16 = 256'h009BFC7E600000000000000003FFFC011C00000000000000C000008000000000;
defparam prom_inst_34.INIT_RAM_17 = 256'h0000000000000060000000000000000000000000000000000000000000000000;
defparam prom_inst_34.INIT_RAM_18 = 256'h000000000000000000000000000000001FF98E7C0000000000000003FFFC000E;
defparam prom_inst_34.INIT_RAM_19 = 256'h723F9F8000000000000001FFFF00238000000000000030000040000000000000;
defparam prom_inst_34.INIT_RAM_1A = 256'h00000000000C0000080000000000000000000000000000000000000000000003;
defparam prom_inst_34.INIT_RAM_1B = 256'h0000000000000000000000000000006CFE1FB000000000000000FFFF9049E000;
defparam prom_inst_34.INIT_RAM_1C = 256'hC7EE000000000000007FFFC087F0000000000000060000000000000000000000;
defparam prom_inst_34.INIT_RAM_1D = 256'h00000001800004000000000000000000000000000000000000000000000009FE;
defparam prom_inst_34.INIT_RAM_1E = 256'h00200000000000000000000000013F1FC7C00000000000003FFFE007FE000000;
defparam prom_inst_34.INIT_RAM_1F = 256'hF80000000000001FFFF008FFC0000000000000C0000080000000000000000000;
defparam prom_inst_34.INIT_RAM_20 = 256'h0000300000800000000000000000000000000000000000000000000000373F8B;
defparam prom_inst_34.INIT_RAM_21 = 256'h00000000000000000000000006FFE1F30000000000000FFFF0087FF800000000;
defparam prom_inst_34.INIT_RAM_22 = 256'h000000000003FFE0003FFF000000000000180000100000000000000000000000;
defparam prom_inst_34.INIT_RAM_23 = 256'h060000000000000000000000000000040000000000000000000000009FC4F3E0;
defparam prom_inst_34.INIT_RAM_24 = 256'h00000000000000000000001B81EC5C000000000001FFE0001FFFA00000000000;
defparam prom_inst_34.INIT_RAM_25 = 256'h000000007FF08007FFF400000000000380000200000000000000000000000000;
defparam prom_inst_34.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000037FF0F98000;
defparam prom_inst_34.INIT_RAM_27 = 256'h000000000000000000006FE3397000000000001FF80000FFFD000000000000C0;
defparam prom_inst_34.INIT_RAM_28 = 256'h00000FFE00003FFF600000000000300000400000000000000000000FC0002000;
defparam prom_inst_34.INIT_RAM_29 = 256'h4000000000000000000004FF0000200000000000000000000009E8FE1E000000;
defparam prom_inst_34.INIT_RAM_2A = 256'h000000000000000001B9F87FC00000000003FF10000FFFC80000000000180000;
defparam prom_inst_34.INIT_RAM_2B = 256'h01FFC00003FFF20000000000060000080000000000000000000E7FF800000000;
defparam prom_inst_34.INIT_RAM_2C = 256'h0000000000000000077FFF8000000000000000000000000017FF8FF000000000;
defparam prom_inst_34.INIT_RAM_2D = 256'h0000000000000006FE23FC000000000063F00008FFF980000000000180000000;
defparam prom_inst_34.INIT_RAM_2E = 256'h7C40007FFE600000000000C00000000000000000000000063FFFF80000000000;
defparam prom_inst_34.INIT_RAM_2F = 256'h00000000000003DFFFFF80000000000000000000000000D88FFF80000000003E;
defparam prom_inst_34.INIT_RAM_30 = 256'h00000000000013BFFFE0000000003B9F00001FFF180000000000300000400000;
defparam prom_inst_34.INIT_RAM_31 = 256'h010FFF8C00000000000C0000000000000000000000013FFFFFF8000000000000;
defparam prom_inst_34.INIT_RAM_32 = 256'h00000000009FFFFFFF800000000000000000000000007FFFF0000000003EFFE1;
defparam prom_inst_34.INIT_RAM_33 = 256'h00000000004FFFFC0000000039BFF81E07FFE700000000000600000000000000;
defparam prom_inst_34.INIT_RAM_34 = 256'hFFF1800000000001800004000000000000000000EFFFFFFFF800000000000000;
defparam prom_inst_34.INIT_RAM_35 = 256'h00000077FFFFFFFF00000000000000000000000004FFFF00000000382FFF8007;
defparam prom_inst_34.INIT_RAM_36 = 256'h00000000FFFF80000000381DFFFD0FFFF8C00000000000200000000000000000;
defparam prom_inst_34.INIT_RAM_37 = 256'h7000000000001800000000000000000000001BFFFFFFFFF00000000000000000;
defparam prom_inst_34.INIT_RAM_38 = 256'h000DFFFFFFFFFF0000000000000000000000000FFFC0000000387EFFFFFFFFF8;
defparam prom_inst_34.INIT_RAM_39 = 256'h000000FFC00000003C3FBFFFFFFFFC3800000000000600000800000000000000;
defparam prom_inst_34.INIT_RAM_3A = 256'h0000000003000002000000000000000006FFFFCFFFFDE0000000000000000000;
defparam prom_inst_34.INIT_RAM_3B = 256'h7FFFE0FFFFBE00000000000000000000000000000000001F1F1FFFFFFFFE3C00;
defparam prom_inst_34.INIT_RAM_3C = 256'h0000000000001FFF07FFFFFFFE1E000000000000C00000000000000000000003;
defparam prom_inst_34.INIT_RAM_3D = 256'h0000003000000000000000000000019FFFF80FFFE7E000000000000000000000;
defparam prom_inst_34.INIT_RAM_3E = 256'hFC00DFFC7E000000000000000000000000000000000FFF01FFFFFFFF0F000000;
defparam prom_inst_34.INIT_RAM_3F = 256'h0000000007FF807FFF7FFF878000000000001C00002000000000000000006FFF;

pROM prom_inst_35 (
    .DO({prom_inst_35_dout_w[30:0],prom_inst_35_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_35.READ_MODE = 1'b1;
defparam prom_inst_35.BIT_WIDTH = 1;
defparam prom_inst_35.RESET_MODE = "SYNC";
defparam prom_inst_35.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_35.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF;
defparam prom_inst_35.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFF;
defparam prom_inst_35.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFF;
defparam prom_inst_35.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFF80000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFC0007C7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFC007C07FFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_11 = 256'hFFFFFFFFFFFC0FC07E007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00FC3E0007FFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_14 = 256'hFFFFFFFE000FFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FF00001FFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_17 = 256'hFFFF00001FC0000FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001FFC000783FFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1A = 256'hF0000FCFC007C03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF800FC0FC07C003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1D = 256'h07C00FC3E0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83F8;
defparam prom_inst_35.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF803F87E000FFE00003FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_20 = 256'h000FF00001FFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003FFE0;
defparam prom_inst_35.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFC0003FF00001FF0000FFFFFFFFFFFFFFFFFC03FFFF;
defparam prom_inst_35.INIT_RAM_23 = 256'hFFF000F9FFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003F80000;
defparam prom_inst_35.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFE00001EF00007C7E007C7FFFFFFFFFFFFFE02007FFFFFF;
defparam prom_inst_35.INIT_RAM_26 = 256'hE07C1FFFFFFFFFFFFFE005E0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001FFF0007C07;
defparam prom_inst_35.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFF8000F87F007E007E3E07FFFFFFFFFFFFF0017C1FFFFFFFFF;
defparam prom_inst_35.INIT_RAM_29 = 256'h01FFFFFFFFFFFFFC079800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800FC03F03F0007FE;
defparam prom_inst_35.INIT_RAM_2B = 256'hFFFFFFFFFFFFCF807E003F3F00007F007FFFFFFFFFFFFF07F0001FFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_2C = 256'hFFFFFFFFFFFFE1F00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0F87E0003FF80000F801F;
defparam prom_inst_35.INIT_RAM_2E = 256'hFFFFFFFFFC0FFF00003F800007E007FFFFFFFFFFFFFC0000007FFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_2F = 256'hFFFFFFFFFF8000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80FF00000E700003C801FFFF;
defparam prom_inst_35.INIT_RAM_31 = 256'hFFFFFFE00F800007FF8003C2007FFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_32 = 256'hFFFFFFFE000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01F00007EFF001E0803FFFFFFF;
defparam prom_inst_35.INIT_RAM_34 = 256'hFFFF007F0003E03F81F0203FFFFFFFFFFFFFFFC000001FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_35 = 256'hFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC019F003F003F8F01819FFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_37 = 256'hF8031F01F0003FF8061C7FFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_38 = 256'hFFC0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00C1F1F80003F801CE1FFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3A = 256'h301FF800007E003E07FFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3B = 256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_35.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF60401FC00003D800F01FFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3D = 256'h3F00001E6003807FFFFFFFFFFFFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3E = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC6180;
defparam prom_inst_35.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF866007F0001E3800C01FFFFFFFFFFFFFFFFF80;

pROM prom_inst_36 (
    .DO({prom_inst_36_dout_w[30:0],prom_inst_36_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_36.READ_MODE = 1'b1;
defparam prom_inst_36.BIT_WIDTH = 1;
defparam prom_inst_36.RESET_MODE = "SYNC";
defparam prom_inst_36.INIT_RAM_00 = 256'h000F0E00F007FFFFFFFFFFFDFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_01 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07C00FF;
defparam prom_inst_36.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC0E0031F0078180E801FFFFFFFFFF0C1FFFFE0000;
defparam prom_inst_36.INIT_RAM_03 = 256'h80206300FFFFFFFFFF80001FFFC000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00C00E1F07;
defparam prom_inst_36.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFC01E0381F3C00870C05FFFFFFFFC000003FFF8000003;
defparam prom_inst_36.INIT_RAM_06 = 256'h383027FFFFFFFE00000007FF0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80740601FC003;
defparam prom_inst_36.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFE00CC1C01E000F80C01FFFFFFFF80000001FFF000000FFF;
defparam prom_inst_36.INIT_RAM_09 = 256'h107FFFFFFF8000000003FE000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC030C70038007C03;
defparam prom_inst_36.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFC0C0CC006001C00C81FFFFFFFC000FE00007FC000003FFFFF;
defparam prom_inst_36.INIT_RAM_0C = 256'hFFFFFFE003FFF0001FF8000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFFFFFC180F001C00B003C07;
defparam prom_inst_36.INIT_RAM_0E = 256'hC0FF00FFFFFF1C601C007007C00E01FFFFFFF803FFFF8001FF000000FFFFFFFF;
defparam prom_inst_36.INIT_RAM_0F = 256'hFFFC03FFFFFC003FE000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01FC03F87FFE1DC01E01C037003007FFF;
defparam prom_inst_36.INIT_RAM_11 = 256'hF00FC0FFF81F007C07018403C01FFFFFFE00FFFFFFC007FC000003FFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_12 = 256'h807FFFFFFC01FF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803;
defparam prom_inst_36.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE00FC03E01FFF03C01BC0E18101900FFFFFFF;
defparam prom_inst_36.INIT_RAM_14 = 256'hF807FFC034023C38C0408407FFFFFFE03FFFFFFF800FF0000007FFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_15 = 256'hFFFFFFF001FE000000E07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF803F81;
defparam prom_inst_36.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFC0700FF87E01FFF00780C3CEE018C107FFFFFFF00F;
defparam prom_inst_36.INIT_RAM_17 = 256'hFFFE01F8303FE00E6043FFFFFFFC07FFFFFFFE007FC000000000FFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_18 = 256'hFFFFC01FF80000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01FC1FE1FC0;
defparam prom_inst_36.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFC03F81F83E0FFFFC0238C03F003E001FFFFFFFE01FFFF;
defparam prom_inst_36.INIT_RAM_1A = 256'hF8083B0038003007FFFFFFFF807FFFFFFFF807FF00000000003FFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_1B = 256'hFE00FFE00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003F03E0707FFF;
defparam prom_inst_36.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFE003C000001FFFFF8307E00E002800FFFFFFFFE03FFFFFFF;
defparam prom_inst_36.INIT_RAM_1D = 256'h407801800E007FFFFFFFF807FFFFFFFFC03FFC00000000007FFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_1E = 256'h0FFF800000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFF8;
defparam prom_inst_36.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFF800000001FFFFFF900700700F803FFFFFFFFF00FFFFFFFFF0;
defparam prom_inst_36.INIT_RAM_20 = 256'hF01C06201FFFFFFFFFC03FFFFFFFFC07FFF00000000000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_21 = 256'hFE00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000007FFFFFF800;
defparam prom_inst_36.INIT_RAM_22 = 256'hFFFFFFFFFFFFF00000003FFFFFFF803F0703041FFFFFFFFFF00FFFFFFFFF01FF;
defparam prom_inst_36.INIT_RAM_23 = 256'hC3810FFFFFFFFFFC00FFFFFFFFC03FFFC00000000007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_24 = 256'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFF80660;
defparam prom_inst_36.INIT_RAM_25 = 256'hFFFFFFFFFFE00000007FFFFFFF0186318047FFFFFFFFFF803FFFFFFFE00FFFF8;
defparam prom_inst_36.INIT_RAM_26 = 256'h13FFFFFFFFFFF00FFFFFFFF007FFFE00000000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_27 = 256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000001FFFFFFFF0606FC0;
defparam prom_inst_36.INIT_RAM_28 = 256'hFFFFFFFFFE000003FFFFFFFF180FE00FFFFFFFFFFFFC01FFFFFFF803FFFF8000;
defparam prom_inst_36.INIT_RAM_29 = 256'hFFFFFFFFFF803FFFFFFE01FFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_2A = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFFFFF300F003FF;
defparam prom_inst_36.INIT_RAM_2B = 256'hFFFFFF8000001FFFFFFFFFC00C00FFFFFFFFFFFFE007FFFFFE00FFFFF8000000;
defparam prom_inst_36.INIT_RAM_2C = 256'hFFFFFFFC01FFFFFF003FFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_2D = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000003FFFFFFFFF003007FFFFF;
defparam prom_inst_36.INIT_RAM_2E = 256'hFFF00000007FFFFFFFFF00C03FFFFFFFFFFFFF803FFFFC001FFFFF8000000000;
defparam prom_inst_36.INIT_RAM_2F = 256'hFFFFE007FFFE000FFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000001FFFFFFFFFE0303FFFFFFFFF;
defparam prom_inst_36.INIT_RAM_31 = 256'h00000003FFFFFFFFFE061FFFFFFFFFFFFFFC01FFF80007FFFFF800000000003F;
defparam prom_inst_36.INIT_RAM_32 = 256'hFF8003CC0003FFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000FFFFFFFFFFE18FFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_34 = 256'h00003FFFFFFFFFFE67FFFFFFFFFFFFFFE000400003FFFFFFC00000000003FFFF;
defparam prom_inst_36.INIT_RAM_35 = 256'h00000007FFFFFFF80000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam prom_inst_36.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_36.INIT_RAM_37 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFF80000007FFFFFFFF00000000007FFFFFFF;
defparam prom_inst_36.INIT_RAM_38 = 256'h000FFFFFFFFFC0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000;
defparam prom_inst_36.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800;
defparam prom_inst_36.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFF80000000007FFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_3B = 256'hFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000003F;
defparam prom_inst_36.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8002F;
defparam prom_inst_36.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFF0000000007FFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_3E = 256'hFFFFFFFE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000001FFFF;
defparam prom_inst_36.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFE0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_37 (
    .DO({prom_inst_37_dout_w[30:0],prom_inst_37_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_37.READ_MODE = 1'b1;
defparam prom_inst_37.BIT_WIDTH = 1;
defparam prom_inst_37.RESET_MODE = "SYNC";
defparam prom_inst_37.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000001FFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_01 = 256'hFFFFF8000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFF;
defparam prom_inst_37.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_04 = 256'hFFF800000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE20007FFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_07 = 256'hFFC0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_08 = 256'hFFFFFFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_0A = 256'h8000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00FFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_0B = 256'hFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFF0000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_0D = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01FFFFFFFFFFFE00;
defparam prom_inst_37.INIT_RAM_0F = 256'hFFFFFFFFFFFFFC007FFFFFFFFFFFC000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_10 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_11 = 256'hFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFC0000;
defparam prom_inst_37.INIT_RAM_12 = 256'hFFFFFFFFE003FFFFFFFFFFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_14 = 256'hFFFFFF801FFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFF0000007;
defparam prom_inst_37.INIT_RAM_15 = 256'hFFF807FFFFFFFFFFFFFFFFFE000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_17 = 256'hFFF0007FFFFFFFFFFFFFFFFFFFFFFFFF003FFFFFFFFFFFFFFFFFFFC000001FFF;
defparam prom_inst_37.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8081FFFFFFF8001FFFFFFFFFFFF8003;
defparam prom_inst_37.INIT_RAM_1A = 256'h0207FFFFFFC0000FFFFFFFFFF003FFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF;
defparam prom_inst_37.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFE000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_37.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE2001FFFFFFE00000FFFFFFFFC0FFFFFFFF;
defparam prom_inst_37.INIT_RAM_1D = 256'h7FFFFFF800000FFFFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFC000001FFFFFFFF;
defparam prom_inst_37.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0080;
defparam prom_inst_37.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC0403FFFFFFC000003FFFFFE0FFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_20 = 256'hFFFF0000007FFFFC1FFFFFFFFFFFFFFFFFFE01FFFFFFFFF0000007FFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_21 = 256'hC0007FFFFFFFFE000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFF;
defparam prom_inst_37.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFC000001FFFF83FFFFFFFFFFF00FFFF;
defparam prom_inst_37.INIT_RAM_23 = 256'hF000000FFFF07FFFFFFFFF8000000000003FFFFFFFFFC000001FFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_24 = 256'hFFFFFFFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFF;
defparam prom_inst_37.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFF0001FFFFFFFC000003FFF0FFFFFFFFF000FFFFFFFFC3;
defparam prom_inst_37.INIT_RAM_26 = 256'h0001FFE1FFFFFFFFC03FFFFFFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_27 = 256'hFFFFFFFFE000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFF80;
defparam prom_inst_37.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFE000FFFFFFFFE00000FFE3FFFFFFFF81FFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_29 = 256'h7FE3FFFFFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFC000001FFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_2A = 256'hFFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFF80000;
defparam prom_inst_37.INIT_RAM_2B = 256'hFFFFFFFFFFFFF8003FFFFFFFFF00003FE3FFFFFFFE0FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_2C = 256'hFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_2D = 256'hFFFE000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFFFFFFFFC0001FE3;
defparam prom_inst_37.INIT_RAM_2E = 256'hFFFFFFFFFF000FFFFFFFFFF8000FE3FFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_2F = 256'hFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_30 = 256'hF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFF000FF3FFFF;
defparam prom_inst_37.INIT_RAM_31 = 256'hFFFFFFC001FFFFFFFFFFC00FF1FFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_32 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_33 = 256'h00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFF80FF9FFFFFFF8;
defparam prom_inst_37.INIT_RAM_34 = 256'hFFF0007FFFFFFFFFFF0FF8FFFFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_37.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_36 = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFCFFFFFFF0FFFF;
defparam prom_inst_37.INIT_RAM_37 = 256'h000FFFFFFFFFFFFFFE7FFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_37.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_37.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFF3FFFFFF0FFFFFFFF;
defparam prom_inst_37.INIT_RAM_3A = 256'hFFFFFFFFFFFFFF9FFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000;
defparam prom_inst_37.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003;
defparam prom_inst_37.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFFFEFFFFFF0FFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_3D = 256'hFFFFFFFFFFF3FFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000003FF;
defparam prom_inst_37.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFF;
defparam prom_inst_37.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFF9FFFFFCFFFFFFFFFFFFFFFF;

pROM prom_inst_38 (
    .DO({prom_inst_38_dout_w[30:0],prom_inst_38_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_38.READ_MODE = 1'b1;
defparam prom_inst_38.BIT_WIDTH = 1;
defparam prom_inst_38.RESET_MODE = "SYNC";
defparam prom_inst_38.INIT_RAM_00 = 256'hFFFFFFFCFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000FFFFF;
defparam prom_inst_38.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFC000001FFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFF;
defparam prom_inst_38.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFE7FFFFE3FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_03 = 256'hFFFF3FFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000003FFFFFFF;
defparam prom_inst_38.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFF0000003FFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFCFFFFF8FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_06 = 256'hE7FFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFFFFFF;
defparam prom_inst_38.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFC000000FFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_08 = 256'hFFFFFFFFFFFFF0003FFFFFFFFFFFFFF3FFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_09 = 256'hFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0A = 256'hFFFFFFFFFFFF0000003FFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFF9FF;
defparam prom_inst_38.INIT_RAM_0B = 256'hFFFFFFFFFC0007FFFFFFFFFFFFFCFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0C = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0D = 256'hFFFFFFFFFC000000FFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFF3FFFFE;
defparam prom_inst_38.INIT_RAM_0E = 256'hFFFFFF0001FFFFFFFFFFFFFF9FFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_10 = 256'hFFFFFFF0000003FFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFCFFFFFCFFF;
defparam prom_inst_38.INIT_RAM_11 = 256'hFFE0003FFFFFFFFFFFFFF7FFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_13 = 256'hFFFFC000000FFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFF9FFFFF3FFFFFF;
defparam prom_inst_38.INIT_RAM_14 = 256'h0007FFFFFFFFFFFFFCFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFFFFFFFFE0078;
defparam prom_inst_38.INIT_RAM_16 = 256'hFF0000001FFFFFFFFFFFFFFFFC00000003FFFFFFFFFFFFFF3FFFFE7FFFFFFFFF;
defparam prom_inst_38.INIT_RAM_17 = 256'hFFFFFFFFFFFFFF9FFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000003FFFFFFFFFFFFFFFC00000001;
defparam prom_inst_38.INIT_RAM_19 = 256'h0000007FFFFFFFFFFFFFFE000000007FFFFFFFFFFFFFCFFFFF9FFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_1A = 256'hFFFFFFFFFFF3FFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_38.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFF000000001FFF;
defparam prom_inst_38.INIT_RAM_1C = 256'h0001FFFFFFFFFFFFFF800000000FFFFFFFFFFFFFF9FFFFF3FFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_1D = 256'hFFFFFFFE7FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam prom_inst_38.INIT_RAM_1E = 256'hFFDFFFFFFFFFFFFFFFFFFFFFFFFE0000003FFFFFFFFFFFFFC000000001FFFFFF;
defparam prom_inst_38.INIT_RAM_1F = 256'h07FFFFFFFFFFFFE0000000003FFFFFFFFFFFFF3FFFFE7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_20 = 256'hFFFFCFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam prom_inst_38.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFF00000000007FFFFFFFF;
defparam prom_inst_38.INIT_RAM_22 = 256'hFFFFFFFFFFFC0000000000FFFFFFFFFFFFE7FFFFCFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_23 = 256'hF9FFFFE7FFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFF0000001F;
defparam prom_inst_38.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFE0000003FFFFFFFFFFFE00000000001FFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_25 = 256'hFFFFFFFF800000000003FFFFFFFFFFFC7FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_26 = 256'hFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFF;
defparam prom_inst_38.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFE00000000000FFFFFFFFFFFF3F;
defparam prom_inst_38.INIT_RAM_28 = 256'hFFFFF000000000001FFFFFFFFFFFCFFFFF3FFFFFFFFFFFFFFFFFFFF03FFFDFFF;
defparam prom_inst_38.INIT_RAM_29 = 256'h9FFFFFFFFFFFFFFFFFFFF800FFFFDFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFF;
defparam prom_inst_38.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFE0000003FFFFFFFFFFC000000000007FFFFFFFFFFE7FFFF;
defparam prom_inst_38.INIT_RAM_2B = 256'hFE000000000001FFFFFFFFFFF9FFFFE7FFFFFFFFFFFFFFFFFFF00007FFFFFFFF;
defparam prom_inst_38.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFFFFFFFE000000FFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFF8000003FFFFFFFFFF8000000000007FFFFFFFFFFE7FFFFBFF;
defparam prom_inst_38.INIT_RAM_2E = 256'h00000000001FFFFFFFFFFF3FFFFCFFFFFFFFFFFFFFFFFFF8000007FFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2F = 256'hFFFFFFFFFFFFFC0000007FFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFC0;
defparam prom_inst_38.INIT_RAM_30 = 256'hFFFFFFFFFFFFE000001FFFFFFFFFC4000000000007FFFFFFFFFFCFFFFF3FFFFF;
defparam prom_inst_38.INIT_RAM_31 = 256'h00000003FFFFFFFFFFF3FFFFDFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_32 = 256'hFFFFFFFFFF000000007FFFFFFFFFFFFFFFFFFFFFFFFE00000FFFFFFFFFC10000;
defparam prom_inst_38.INIT_RAM_33 = 256'hFFFFFFFFFF800003FFFFFFFFC6400000000000FFFFFFFFFFF9FFFFF7FFFFFFFF;
defparam prom_inst_38.INIT_RAM_34 = 256'h00007FFFFFFFFFFE7FFFF9FFFFFFFFFFFFFFFFFF0000000007FFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_35 = 256'hFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFF80000FFFFFFFFC7D0000000;
defparam prom_inst_38.INIT_RAM_36 = 256'hFFFFFFFF00007FFFFFFFC7E200000000003FFFFFFFFFFF9FFFFE7FFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_37 = 256'h0FFFFFFFFFFFE7FFFF9FFFFFFFFFFFFFFFFFE0000000000FFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_38 = 256'hFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFC7810000000000;
defparam prom_inst_38.INIT_RAM_39 = 256'hFFFFFF003FFFFFFFC3C0400000000007FFFFFFFFFFF9FFFFE7FFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3A = 256'hFFFFFFFFFCFFFFF9FFFFFFFFFFFFFFFFF800000000001FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3B = 256'h000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0E0000000000003FF;
defparam prom_inst_38.INIT_RAM_3C = 256'hFFFFFFFFFFFFE000000000000001FFFFFFFFFFFF3FFFFEFFFFFFFFFFFFFFFFFC;
defparam prom_inst_38.INIT_RAM_3D = 256'hFFFFFFCFFFFFBFFFFFFFFFFFFFFFFE0000000000001FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3E = 256'h0000200001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000FFFFFF;
defparam prom_inst_38.INIT_RAM_3F = 256'hFFFFFFFFF8000000000000007FFFFFFFFFFFE3FFFFCFFFFFFFFFFFFFFFFF8000;

pROM prom_inst_39 (
    .DO({prom_inst_39_dout_w[30:0],prom_inst_39_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_39.READ_MODE = 1'b1;
defparam prom_inst_39.BIT_WIDTH = 1;
defparam prom_inst_39.RESET_MODE = "SYNC";
defparam prom_inst_39.INIT_RAM_00 = 256'hFE0080000F0008BC35C000001F2F6FFDFCF5D8F1A7FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_01 = 256'h7F3C3F197FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FF543A81BB905E5C0007FFFB;
defparam prom_inst_39.INIT_RAM_02 = 256'hFFFFC9FF8FD5F0E7EC16AE000087FF0E03800001C0000D0D0000000F9537FFFF;
defparam prom_inst_39.INIT_RAM_03 = 256'h900001F000000C18000007C2BFFFFFBFF3CBFD6FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_04 = 256'h7DAB207FFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFE7FCBF58F80D5B800423FE3F80;
defparam prom_inst_39.INIT_RAM_05 = 256'hF05FE4FFE3AC43C354C00000F919E00C00003800005300000003F237FFFFDFEF;
defparam prom_inst_39.INIT_RAM_06 = 256'h001E00000000000000F8537FFFE7F7F79B3A27FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_07 = 256'hD7717FFFFFFFFFFFFFFFFFFFFFFFFFF82BED6BF26E2203D570000267D8600100;
defparam prom_inst_39.INIT_RAM_08 = 256'h3130DE292407B558000000020006400005800002000000007CDA7DF7FBFBFEFF;
defparam prom_inst_39.INIT_RAM_09 = 256'hE00000000000001F28B71FFDFCFEFFF2037FFFFFFFFFFFFFFFFFFFFFFFFFFC07;
defparam prom_inst_39.INIT_RAM_0A = 256'h31FFFFFFFFFFFFFFFFFFFFFFFFFF07E27E83009380FDD7000000008001500003;
defparam prom_inst_39.INIT_RAM_0B = 256'hC0644E8C2F75C0000182000074000078000000000000079B7FF6FEFF7F7E7D2D;
defparam prom_inst_39.INIT_RAM_0C = 256'h000000000003C5CFF5FFBFBF9FB792069FFFFFFFFFFFFFFFFFFFFFFFFC01FC1F;
defparam prom_inst_39.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFE1003F9FC00105A007DF6000000000001700003E00;
defparam prom_inst_39.INIT_RAM_0E = 256'h11F903F7D8000000000000C0000F00000000000000F17BFFFFDFDFEFFF7DFC05;
defparam prom_inst_39.INIT_RAM_0F = 256'h000000007C19FFEFEFF7F7EFEFB4EC1FBFFFFFFFFFFFFFFFFFFFFD202FF3E000;
defparam prom_inst_39.INIT_RAM_10 = 256'hBFFFFFFFFFFFFFFFFFFC500FFA3000041900FD26000000000000700007C00000;
defparam prom_inst_39.INIT_RAM_11 = 256'hA01E498000000000000C0001F00000000000003F487FF33BFBFBFFFFFF0A53FC;
defparam prom_inst_39.INIT_RAM_12 = 256'h000007923F8DFCFDFEFDFDFFD48E33FFFFFFDFFFFFFFFFFFFF5401FE00C3C1F8;
defparam prom_inst_39.INIT_RAM_13 = 256'hFFEEFFFFFFFFFFFEC400FFC00000BE000192600000000000320000DC00000000;
defparam prom_inst_39.INIT_RAM_14 = 256'h6C9800000000000980003700000000000003E4C7D32B9F7F7FFFFFFE0F50F357;
defparam prom_inst_39.INIT_RAM_15 = 256'h00F978E482B9FFBFD3EDFFF238100FFFFF9FFFFFFFFFFFB0002FE00000078000;
defparam prom_inst_39.INIT_RAM_16 = 256'h99FFFFFFFFFD1C000EF800000060000BEC000000000000E00017C00000000000;
defparam prom_inst_39.INIT_RAM_17 = 256'h000000000000BC0007600000000000003E4FD0C60BDFEFD0A0B7FEA78F03FFFF;
defparam prom_inst_39.INIT_RAM_18 = 256'h91FAEFE126F7F0180A7FC772C0393FFDDFFFFFFFF6772001FC000000000003FB;
defparam prom_inst_39.INIT_RAM_19 = 256'hFFFFFFFFFAC0005F000000000001E4C000000000000E0001B80000000000000F;
defparam prom_inst_39.INIT_RAM_1A = 256'h00000000178000AE00000000000001E67F9002105FF8040017FC54E0000DEEFB;
defparam prom_inst_39.INIT_RAM_1B = 256'hD60039847E020000BFF7FA00007DBCFF7FF7FF63080013E000000000005D6000;
defparam prom_inst_39.INIT_RAM_1C = 256'hF7B77F200002F0000000000037D8000000000000E0003B80000000000000798F;
defparam prom_inst_39.INIT_RAM_1D = 256'h00000178001DC00000000000001F63FD0001940E01000047FDE380003BA7BBDF;
defparam prom_inst_39.INIT_RAM_1E = 256'h000D43C0400001EF3C5C000277F0BFFFFC58180800DF00000000015FAC000000;
defparam prom_inst_39.INIT_RAM_1F = 256'h58A6880011E0000000006F930000000000005E00053000000000000003CCFF95;
defparam prom_inst_39.INIT_RAM_20 = 256'h0027C0039C00000000000001FB17DAD000D6E82000007BFDFAA0003E9E8FADD5;
defparam prom_inst_39.INIT_RAM_21 = 256'h01729000001DBFFF62000637A1239DA2008000077E1000000061D58000000000;
defparam prom_inst_39.INIT_RAM_22 = 256'h000000E3E7000000BDFAE0000000000009E000B7000000000000007E23FF4D30;
defparam prom_inst_39.INIT_RAM_23 = 256'hB8007B8000000000000007CCB7D79F839824000007F40FEB30001054A7274022;
defparam prom_inst_39.INIT_RAM_24 = 256'hA0000001FAB03FE600001809C50110C000003C7CFD4001F8FD70000000000004;
defparam prom_inst_39.INIT_RAM_25 = 256'h0003D7DD408AB47A98000000000001FE001EE000000000000001F99A3F70E781;
defparam prom_inst_39.INIT_RAM_26 = 256'h15B0000000000000003E3287DD6046BE000000FDFBE71EE00000008801800000;
defparam prom_inst_39.INIT_RAM_27 = 256'h000032FFFED79C00000848000000000000F93EB9E3CC8D4E00000000000173C0;
defparam prom_inst_39.INIT_RAM_28 = 256'h0F93F81AC9C6AF0000000000007CF00FDC000000000000000FE77B359C007960;
defparam prom_inst_39.INIT_RAM_29 = 256'h8000000000000001F869B3F9E1015600000FFFFFBAF180000008040040000000;
defparam prom_inst_39.INIT_RAM_2A = 256'h0ADFFFEE9A2000000000000000000001F98FF00D77B78000000000003FBE03E7;
defparam prom_inst_39.INIT_RAM_2B = 256'h88800956B38000000000001AE781EDC0000000000000003F0ED5FB96BBF7A000;
defparam prom_inst_39.INIT_RAM_2C = 256'h0000000000000FF0CACFBB773EFA0001E7FFFAADC6000000000000000000001F;
defparam prom_inst_39.INIT_RAM_2D = 256'hFFFFA3F08000000000000000000003F89016EEB3C000000000000F3DFFFC6000;
defparam prom_inst_39.INIT_RAM_2E = 256'hBE1F33C0000000000007DA7DFFBC0000000000000000FE1C83FBA7FFF38000D9;
defparam prom_inst_39.INIT_RAM_2F = 256'h00000000001FE18CFFB93FD050006CFFFF7AFEB0000000000000000000003F86;
defparam prom_inst_39.INIT_RAM_30 = 256'hFEF6240000000000000000000001FC1C21C3E0000000000001C39FFECF000000;
defparam prom_inst_39.INIT_RAM_31 = 256'h0FE0000000000000736FFE91C00000000000000007FE19F7FD73C89040373FFF;
defparam prom_inst_39.INIT_RAM_32 = 256'h00000000FFE39C5F962417207B8FFFEBBFC000000000000000000000001FF000;
defparam prom_inst_39.INIT_RAM_33 = 256'hF8E80000000000000000000000FFFEFFE00000000000003BD3FF807000000000;
defparam prom_inst_39.INIT_RAM_34 = 256'h0000000000001FFCFFC0BC00000000000000000FFC39FDFB14376A8EC3FFF4EF;
defparam prom_inst_39.INIT_RAM_35 = 256'h000000FFC399FFF680767FE0FFFD7A3EBC00000000000000000000000FFFFF80;
defparam prom_inst_39.INIT_RAM_36 = 256'hC000000000000000000000007FFF8000000000000007BA7FF42F000000000000;
defparam prom_inst_39.INIT_RAM_37 = 256'h0000000002FE1FFC3BC000000000000000003FFE3BBDBCDC0C99F01FFEFF92AF;
defparam prom_inst_39.INIT_RAM_38 = 256'h0003FFE31FD0E782873C07FFAF7F1AC000000000000000000000000000000000;
defparam prom_inst_39.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000FD8FFE00F000000000000000;
defparam prom_inst_39.INIT_RAM_3A = 256'h0000001F87FFC33C0000000000000000007FFE33FC0EB85FDE41FFD9DFE93A00;
defparam prom_inst_39.INIT_RAM_3B = 256'h07FFE31FC06ACB7AC0FFF67FFE26400000000000000000000000000000000000;
defparam prom_inst_39.INIT_RAM_3C = 256'h00000000000000000000000000000000000003FFFFE9DE000000000000000000;
defparam prom_inst_39.INIT_RAM_3D = 256'h00007FFFF877C00000000000000000007FFF39500EA0E6583FFD3AFFE3900000;
defparam prom_inst_39.INIT_RAM_3E = 256'hFFF19C00EF50DB0FFF5CFFFC3400000000000000000000000000000000000000;
defparam prom_inst_39.INIT_RAM_3F = 256'h000000000000000000000000000000000007F17E11C000000000000000000017;

pROM prom_inst_40 (
    .DO({prom_inst_40_dout_w[30:0],prom_inst_40_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_40.READ_MODE = 1'b1;
defparam prom_inst_40.BIT_WIDTH = 1;
defparam prom_inst_40.RESET_MODE = "SYNC";
defparam prom_inst_40.INIT_RAM_00 = 256'hFFF87FFFF8FFFFFFFFFFFFFFE011FFFE0011FF09FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_01 = 256'h017EC09DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000A617E646F85C3FFFFFFFF;
defparam prom_inst_40.INIT_RAM_02 = 256'hFFFFFE00103C0F1813E061FFFFFFFFFFFD3FFFFF3FFFFFFFFFFFFFF01CFFFF00;
defparam prom_inst_40.INIT_RAM_03 = 256'h2FFFFE4FFFFFFFFFFFFFF80D7FFF800017E41DDFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_04 = 256'h7F47EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00180380A387F0B87FFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_05 = 256'hFFA00B801853BCFC2C3FFFFFFFFFFFCBFFFF87FFFFFFFFFFFFFC019FFFC00001;
defparam prom_inst_40.INIT_RAM_06 = 256'hFFE1FFFFFFFFFFFFFF008FFFF0000017F4FDFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_07 = 256'h7F8BFFFFFFFFFFFFFFFFFFFFFFFFFFFFD40A940CC1DDF40B0FFFFFFFFFFFF8FF;
defparam prom_inst_40.INIT_RAM_08 = 256'h8687E1FC9BFC42C7FFFFFFFFFFFA3FFFFA7FFFFFFFFFFFFF80BFBDF00000017F;
defparam prom_inst_40.INIT_RAM_09 = 256'h1FFFFFFFFFFFFFE03F7F1E00000017F9FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_40.INIT_RAM_0A = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFFFA11C182FE7C7F0030FFFFFFFFFFFE0FFFFC;
defparam prom_inst_40.INIT_RAM_0B = 256'h407BB973D00C3FFFFFFFFFFFA3FFFF07FFFFFFFFFFFFF817FF7700000000FF91;
defparam prom_inst_40.INIT_RAM_0C = 256'hFFFFFFFFFFFC07FFFD800000007FF11BFFFFFFFFFFFFFFFFFFFFFFFFFFFE03C0;
defparam prom_inst_40.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF80600001FA5FF0031FFFFFFFFFFFE4FFFFE1FF;
defparam prom_inst_40.INIT_RAM_0E = 256'h1A06FE00C7FFFFFFFFFFF83FFFF4FFFFFFFFFFFFFF03FFFF600000001FFF21F7;
defparam prom_inst_40.INIT_RAM_0F = 256'hFFFFFFFF80DFFFF40000001FFFFC37FFFFFFFFFFFFFFFFFFFFFFFFFFC00E0000;
defparam prom_inst_40.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFF405E0000026FF80E1FFFFFFFFFFFF0FFFF93FFFFF;
defparam prom_inst_40.INIT_RAM_11 = 256'h5FF0387FFFFFFFFFFF83FFFE0FFFFFFFFFFFFFC05FFFF780000007FFFFC3FFFF;
defparam prom_inst_40.INIT_RAM_12 = 256'hFFFFF817FF8EFA000003FFFFFC3EFFFFFFFFFFFFFFFFFFFFFFFFFD01FFFFC003;
defparam prom_inst_40.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFF403FFFFF81FFFE261FFFFFFFFFFFD1FFFF23FFFFFFFF;
defparam prom_inst_40.INIT_RAM_14 = 256'hC187FFFFFFFFFFF27FFFC8FFFFFFFFFFFFFC075FD3BBE00001FFFFFE846FFFFF;
defparam prom_inst_40.INIT_RAM_15 = 256'hFF0187E4C3BC000053EDFFFA47E7FFFFFFFFFFFFFFFFFFFFFFC01FFFFFFCFFFF;
defparam prom_inst_40.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFF107FFFFFFDFFFF863FFFFFFFFFFFC1FFFE83FFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_17 = 256'hFFFFFFFFFFFF03FFF81FFFFFFFFFFFFFC07030F71BC00030A0B7FFE079FFFFFF;
defparam prom_inst_40.INIT_RAM_18 = 256'h1E06FFE1A50010180A7FFD857FFFFFFFFFFFFFFFFFFFFFFF83FFFFFFFFFFFD18;
defparam prom_inst_40.INIT_RAM_19 = 256'hFFFFFFFFFFFFFF80FFFFFFFFFFFE0C3FFFFFFFFFFFC1FFFE47FFFFFFFFFFFFF0;
defparam prom_inst_40.INIT_RAM_1A = 256'hFFFFFFFFE07FFF41FFFFFFFFFFFFFE07815FFE187000040017FF681FFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1B = 256'h2FFFF98602020000BF0903FFFFFFFFFFFFFFFFFFFFFFEC1FFFFFFFFFFFA31FFF;
defparam prom_inst_40.INIT_RAM_1C = 256'hFFFFFFFFFFFC0FFFFFFFFFFDCAC7FFFFFFFFFFF81FFFC07FFFFFFFFFFFFF81F0;
defparam prom_inst_40.INIT_RAM_1D = 256'hFFFFFE07FFE23FFFFFFFFFFFFFE07C03DFFF9C2001000047C0586FFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1E = 256'hFFFDC2C0400001E00393FFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFE463FFFFFF;
defparam prom_inst_40.INIT_RAM_1F = 256'hFFFFFFFFE21FFFFFFFFF7030FFFFFFFFFFFFC1FFF80FFFFFFFFFFFFFFC0F007F;
defparam prom_inst_40.INIT_RAM_20 = 256'hFFC83FFC43FFFFFFFFFFFFFE03E227FFFFDEF82000007C00155FFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_21 = 256'hFFF39000001E40009DFFFFFFFFFFFFFFFFFFFFF8C1FFFFFFFFF02C7FFFFFFFFF;
defparam prom_inst_40.INIT_RAM_22 = 256'hFFFFFF041EFFFFFFE0061FFFFFFFFFFFF81FFF10FFFFFFFFFFFFFF803CE4DB3F;
defparam prom_inst_40.INIT_RAM_23 = 256'h07FF907FFFFFFFFFFFFFF80F006FFFFE7C3C0000079BF007CFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_24 = 256'hE0000001CF7FC1F9FFFFFFFFFFFFFFFFFFFFC102EFFFFF78030FFFFFFFFFFFF8;
defparam prom_inst_40.INIT_RAM_25 = 256'hFFFC00355FFFB80587FFFFFFFFFFFE81FFE21FFFFFFFFFFFFFFE01E0AEBEF00F;
defparam prom_inst_40.INIT_RAM_26 = 256'hEA8FFFFFFFFFFFFFFFC03D68E390007E000000F3FFF87F1FFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_27 = 256'h00003DFFFF1FE7FFFFFFFFFFFFFFFFFFFF0041BCFFF012C1FFFFFFFFFFFE803F;
defparam prom_inst_40.INIT_RAM_28 = 256'hF0100787F09860FFFFFFFFFFFF800FF003FFFFFFFFFFFFFFF00782CE7F000760;
defparam prom_inst_40.INIT_RAM_29 = 256'h7FFFFFFFFFFFFFFE007040676000B200000E7FFFC3FEFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2A = 256'h0A3FFFF0FFCFFFFFFFFFFFFFFFFFFFFE01100FF099707FFFFFFFFFFFC081FC50;
defparam prom_inst_40.INIT_RAM_2B = 256'h08FFF039707FFFFFFFFFFFE0207E143FFFFFFFFFFFFFFFC00F4406740009E000;
defparam prom_inst_40.INIT_RAM_2C = 256'hFFFFFFFFFFFFF000F0306740C09E00019FFFFC1FF9FFFFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_40.INIT_RAM_2D = 256'hFFFE07FD7FFFFFFFFFFFFFFFFFFFFC00D021F0703FFFFFFFFFFFF01C000A1FFF;
defparam prom_inst_40.INIT_RAM_2E = 256'h3FE4F03FFFFFFFFFFFF806020083FFFFFFFFFFFFFFFF001F0E06740041C000E7;
defparam prom_inst_40.INIT_RAM_2F = 256'hFFFFFFFFFFE001F0806440203C0063FFFF83FF0FFFFFFFFFFFFFFFFFFFFFC007;
defparam prom_inst_40.INIT_RAM_30 = 256'hC0FFC3FFFFFFFFFFFFFFFFFFFFFE001FDFC01FFFFFFFFFFFFE01800220FFFFFF;
defparam prom_inst_40.INIT_RAM_31 = 256'h001FFFFFFFFFFFFF8CE000883FFFFFFFFFFFFFFFF8001E0002E43066C038FFFF;
defparam prom_inst_40.INIT_RAM_32 = 256'hFFFFFFFF0003E1806E5820387C7FFFF03FF2BFFFFFFFFFFFFFFFFFFFFFE00000;
defparam prom_inst_40.INIT_RAM_33 = 256'hFCD7FFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFFC03000060FFFFFFFFF;
defparam prom_inst_40.INIT_RAM_34 = 256'hFFFFFFFFFFFFE10C000183FFFFFFFFFFFFFFFFF0003E2004BA00078E3FFFF80F;
defparam prom_inst_40.INIT_RAM_35 = 256'hFFFFFF0003E6000F08005F1FFFFE01FF3BFFFFFFFFFFFFFFFFFFFFFFF000007F;
defparam prom_inst_40.INIT_RAM_36 = 256'h7FFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFF846000420FFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_37 = 256'hFFFFFFFFFD010001083FFFFFFFFFFFFFFFFFC0003C4043E0005F8FFFFF00FFCF;
defparam prom_inst_40.INIT_RAM_38 = 256'hFFFC0003E00F540009C3FFFFC07FF6EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0180004C0FFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3A = 256'hFFFFFFE000001303FFFFFFFFFFFFFFFFFF80003C01F1A00021FFFFE00FFCBDFF;
defparam prom_inst_40.INIT_RAM_3B = 256'hF80003E03F9A00063FFFF807FFE7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000008C1FFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3D = 256'hFFFF800002103FFFFFFFFFFFFFFFFFFF80003E13F1B00087FFFE01FFFCFFFFFF;
defparam prom_inst_40.INIT_RAM_3E = 256'h0001E03F1E0010FFFF81FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80E80883FFFFFFFFFFFFFFFFFFFE8;

pROM prom_inst_41 (
    .DO({prom_inst_41_dout_w[30:0],prom_inst_41_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_41.READ_MODE = 1'b1;
defparam prom_inst_41.BIT_WIDTH = 1;
defparam prom_inst_41.RESET_MODE = "SYNC";
defparam prom_inst_41.INIT_RAM_00 = 256'h0006000000000000000000000037FFFE000DFF07E00000000000000000000000;
defparam prom_inst_41.INIT_RAM_01 = 256'h00FEC07C00000000000000000000000000000003FFE19FFF9FFFE3C000000000;
defparam prom_inst_41.INIT_RAM_02 = 256'h000001FFE003FFE7FFF9E000000000000080000000000000000000000BFFFF00;
defparam prom_inst_41.INIT_RAM_03 = 256'h60000040000000000000000EFFFF80000FE803C0000000000000000000000000;
defparam prom_inst_41.INIT_RAM_04 = 256'hFF801C000000000000000000000000000000FFE0007FFC7DFE78000000000000;
defparam prom_inst_41.INIT_RAM_05 = 256'h005FF00027FC033F9C0000000000001800000000000000000000037FFFE00000;
defparam prom_inst_41.INIT_RAM_06 = 256'h00100000000000000001FFFFF000000FF800C000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_07 = 256'h8018000000000000000000000000000003F060033E000FE70000000000000C00;
defparam prom_inst_41.INIT_RAM_08 = 256'h78780013C003F9C00000000000010000000000000000000000E1FDF0000000FF;
defparam prom_inst_41.INIT_RAM_09 = 256'h800000000000000010FF1C0000000FFC03800000000000000000000000000008;
defparam prom_inst_41.INIT_RAM_0A = 256'h7800000000000000000000000000000C3E7C018000FE70000000000000C00000;
defparam prom_inst_41.INIT_RAM_0B = 256'hBF8000003F9C00000000000010000000000000000000001C3FF700000001FFC2;
defparam prom_inst_41.INIT_RAM_0C = 256'h000000000000021FFD800000007FFCE78000000000000000000000000001003F;
defparam prom_inst_41.INIT_RAM_0D = 256'h00000000000000000000000000401FFFFE00000FE70000000000000C00000000;
defparam prom_inst_41.INIT_RAM_0E = 256'hE40001F9C0000000000002000000000000000000000287FFC00000003FFF9E70;
defparam prom_inst_41.INIT_RAM_0F = 256'h0000000000E3FFF80000000FFFFBC7000000000000000000000000001001FFFF;
defparam prom_inst_41.INIT_RAM_10 = 256'h000000000000000000000000001FFFFFC0007E60000000000001800001000000;
defparam prom_inst_41.INIT_RAM_11 = 256'h000F98000000000000600001000000000000000070FFF7C0000007FFFFBC7000;
defparam prom_inst_41.INIT_RAM_12 = 256'h0000001C7F8FFC000003FFFFFBC6000000000000000000000000000000003FFC;
defparam prom_inst_41.INIT_RAM_13 = 256'h00000000000000000000000000007E0001CE0000000000000800000000000000;
defparam prom_inst_41.INIT_RAM_14 = 256'h33800000000000060000080000000000000007BFD3BBC00000FFFFFEF8E00000;
defparam prom_inst_41.INIT_RAM_15 = 256'h0001FFE4C3BE000053EDFFFD8E1C000000000000000000000010000000030000;
defparam prom_inst_41.INIT_RAM_16 = 256'h00000000000000000400000000000004E0000000000001000008000000000000;
defparam prom_inst_41.INIT_RAM_17 = 256'h000000000000C0000000000000000000007FF0F71BE00030A0B7FFD8E8000000;
defparam prom_inst_41.INIT_RAM_18 = 256'h1FFEFFE1A60000180A7FFE084000000000000000000000010000000000000038;
defparam prom_inst_41.INIT_RAM_19 = 256'h00000000000000200000000000001C0000000000003000004000000000000000;
defparam prom_inst_41.INIT_RAM_1A = 256'h000000000C0000400000000000000007FFDFFE186000040017FCF00000000000;
defparam prom_inst_41.INIT_RAM_1B = 256'hFFFFF98702020000BF0786000000000000000000000008000000000000070000;
defparam prom_inst_41.INIT_RAM_1C = 256'h00000000000100000000000201C00000000000020000000000000000000001FF;
defparam prom_inst_41.INIT_RAM_1D = 256'h00000180000200000000000000007FFFDFFF9C3101000047C03C600000000000;
defparam prom_inst_41.INIT_RAM_1E = 256'hFFFDC340400001F001EF0000000000000000000000200000000000C0E0000000;
defparam prom_inst_41.INIT_RAM_1F = 256'h00000000040000000001907000000000000020000200000000000000000FFFFF;
defparam prom_inst_41.INIT_RAM_20 = 256'h00180000000000000000000003F9FFFFFFDEF820000078000FF0000000000000;
defparam prom_inst_41.INIT_RAM_21 = 256'hFFF39000001E00007F00000000000000000000008000000000281C0000000000;
defparam prom_inst_41.INIT_RAM_22 = 256'h0000000803000000780E0000000000000C00001000000000000000003E1FDF3F;
defparam prom_inst_41.INIT_RAM_23 = 256'h00000000000000000000000FC9FFFFFC7C3C00000700000FE000000000000000;
defparam prom_inst_41.INIT_RAM_24 = 256'hE0000001C00001FE000000000000000000000181B68000D00700000000000003;
defparam prom_inst_41.INIT_RAM_25 = 256'h0000180FE085D00380000000000000400000000000000000000001F11FFEF807;
defparam prom_inst_41.INIT_RAM_26 = 256'h028000000000000000003E07FFE0007E000000E000007FC00000000000000000;
defparam prom_inst_41.INIT_RAM_27 = 256'h00003800000FFC00000000000000000000018043B92001C00000000000008800;
defparam prom_inst_41.INIT_RAM_28 = 256'h001C007C0001E000000000000002000000000000000000000007C43FF8000760;
defparam prom_inst_41.INIT_RAM_29 = 256'h0000000000000000007C27FF80007600000C000003FF80000000000000000000;
defparam prom_inst_41.INIT_RAM_2A = 256'h0B000000FFE00000000000000000000001E0000000F000000000000000800050;
defparam prom_inst_41.INIT_RAM_2B = 256'h0F000000F0000000000000002000040000000000000000000FB2FFF80007E000;
defparam prom_inst_41.INIT_RAM_2C = 256'h0000000000000000FC6FFF80003E00018000003FFC0000000000000000000000;
defparam prom_inst_41.INIT_RAM_2D = 256'h00000FFF800000000000000000000000EFC001F0000000000000010C000A0000;
defparam prom_inst_41.INIT_RAM_2E = 256'hC003F000000000000000060000800000000000000000001FF1FFF80003C000C0;
defparam prom_inst_41.INIT_RAM_2F = 256'h00000000000001FF7FFD80003C0070000001FFF0000000000000000000000007;
defparam prom_inst_41.INIT_RAM_30 = 256'h007FFE0000000000000000000000001FFFC00000000000000001800220000000;
defparam prom_inst_41.INIT_RAM_31 = 256'h000000000000000008600008000000000000000000001FFFFFF80002C0380000;
defparam prom_inst_41.INIT_RAM_32 = 256'h000000000003FEFFFF8000787C0000001FFF8000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_33 = 256'hFFF0000000000000000000000000000000000000000000003000020000000000;
defparam prom_inst_41.INIT_RAM_34 = 256'h000000000000010C000080000000000000000000003FDFFFA000078E00000007;
defparam prom_inst_41.INIT_RAM_35 = 256'h0000000003F9FFFC0000FF00000003FFFE000000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_36 = 256'hC000000000000000000000000000000000000000000002000460000000000000;
defparam prom_inst_41.INIT_RAM_37 = 256'h00000000000100011800000000000000000000003FBFFFC0000F80000000FFFF;
defparam prom_inst_41.INIT_RAM_38 = 256'h00000003FFFFF70001C00000003FFEF000000000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000018000440000000000000000;
defparam prom_inst_41.INIT_RAM_3A = 256'h000000000000010000000000000000000000003FFFFFB000300000001FFEBE00;
defparam prom_inst_41.INIT_RAM_3B = 256'h000003FFFFFB000400000007FFCF800000000000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000840000000000000000000;
defparam prom_inst_41.INIT_RAM_3D = 256'h0000000002300000000000000000000000003FEFFFA00080000003FFFE700000;
defparam prom_inst_41.INIT_RAM_3E = 256'h0001FFFFFE0030000000FFFFEC00000000000000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000080000000000000000000000;

pROM prom_inst_42 (
    .DO({prom_inst_42_dout_w[30:0],prom_inst_42_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_42.READ_MODE = 1'b1;
defparam prom_inst_42.BIT_WIDTH = 1;
defparam prom_inst_42.RESET_MODE = "SYNC";
defparam prom_inst_42.INIT_RAM_00 = 256'hFFF9FFFFF3FFFFFFFFFFFFFFFFC00000000200001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_01 = 256'h00010003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000003FFFFFFFFF;
defparam prom_inst_42.INIT_RAM_02 = 256'hFFFFFE000000000000001FFFFFFFFFFFFE7FFFFCFFFFFFFFFFFFFFFFE0000000;
defparam prom_inst_42.INIT_RAM_03 = 256'h9FFFFF3FFFFFFFFFFFFFFFF0000000000010003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_04 = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_05 = 256'hFF8000000000000003FFFFFFFFFFFFE7FFFFDFFFFFFFFFFFFFFFFC0000000000;
defparam prom_inst_42.INIT_RAM_06 = 256'hFFE7FFFFFFFFFFFFFFFE00000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_07 = 256'h0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFF3FF;
defparam prom_inst_42.INIT_RAM_08 = 256'h000000000000003FFFFFFFFFFFFCFFFFF9FFFFFFFFFFFFFFFF00020800000000;
defparam prom_inst_42.INIT_RAM_09 = 256'h7FFFFFFFFFFFFFFFC000E00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_42.INIT_RAM_0A = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFF3FFFFE;
defparam prom_inst_42.INIT_RAM_0B = 256'h000000000003FFFFFFFFFFFFCFFFFFBFFFFFFFFFFFFFFFE00008000000000000;
defparam prom_inst_42.INIT_RAM_0C = 256'hFFFFFFFFFFFFF80002000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFE0000;
defparam prom_inst_42.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFF3FFFFCFFF;
defparam prom_inst_42.INIT_RAM_0E = 256'h000000003FFFFFFFFFFFFDFFFFF3FFFFFFFFFFFFFFFC0000000000000000000F;
defparam prom_inst_42.INIT_RAM_0F = 256'hFFFFFFFFFF00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000;
defparam prom_inst_42.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFE7FFFFCFFFFFF;
defparam prom_inst_42.INIT_RAM_11 = 256'h000007FFFFFFFFFFFF9FFFFE7FFFFFFFFFFFFFFF800008000000000000000FFF;
defparam prom_inst_42.INIT_RAM_12 = 256'hFFFFFFE000700000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFE0000000000;
defparam prom_inst_42.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFE7FFFF9FFFFFFFFF;
defparam prom_inst_42.INIT_RAM_14 = 256'h007FFFFFFFFFFFF9FFFFE7FFFFFFFFFFFFFFF8002C44000000000001001FFFFF;
defparam prom_inst_42.INIT_RAM_15 = 256'hFFFE001B3C4000002C12000001E3FFFFFFFFFFFFFFFFFFFFFFE0000000000000;
defparam prom_inst_42.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFEFFFFF3FFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_17 = 256'hFFFFFFFFFFFF3FFFFCFFFFFFFFFFFFFFFF800F08E400000F5F48000010FFFFFF;
defparam prom_inst_42.INIT_RAM_18 = 256'hE001001E58000FE7F58000003FFFFFFFFFFFFFFFFFFFFFFE0000000000000007;
defparam prom_inst_42.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFCFFFFF3FFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1A = 256'hFFFFFFFFF3FFFF9FFFFFFFFFFFFFFFF8002001E78007FBFFE800001FFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1B = 256'h0000067801FDFFFF400001FFFFFFFFFFFFFFFFFFFFFFF000000000000000FFFF;
defparam prom_inst_42.INIT_RAM_1C = 256'hFFFFFFFFFFFE000000000000003FFFFFFFFFFFFDFFFFE7FFFFFFFFFFFFFFFE00;
defparam prom_inst_42.INIT_RAM_1D = 256'hFFFFFE7FFFF9FFFFFFFFFFFFFFFF8000200063C0FEFFFFB800001FFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1E = 256'h00023C3FBFFFFE000000FFFFFFFFFFFFFFFFFFFFFFC00000000000001FFFFFFF;
defparam prom_inst_42.INIT_RAM_1F = 256'hFFFFFFFFF80000000000000FFFFFFFFFFFFF9FFFFCFFFFFFFFFFFFFFFFF00000;
defparam prom_inst_42.INIT_RAM_20 = 256'hFFE7FFFF3FFFFFFFFFFFFFFFFC000000002107DFFFFF8000000FFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_21 = 256'h000C6FFFFFE0000000FFFFFFFFFFFFFFFFFFFFFF00000000000003FFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_22 = 256'hFFFFFFF0000000000001FFFFFFFFFFFFF3FFFFCFFFFFFFFFFFFFFFFFC00020C0;
defparam prom_inst_42.INIT_RAM_23 = 256'hFFFFE7FFFFFFFFFFFFFFFFF00000000003C3FFFFF80000001FFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_24 = 256'h1FFFFFFE00000001FFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFC;
defparam prom_inst_42.INIT_RAM_25 = 256'hFFFFE000000000007FFFFFFFFFFFFF3FFFF9FFFFFFFFFFFFFFFFFE0000010000;
defparam prom_inst_42.INIT_RAM_26 = 256'hFC7FFFFFFFFFFFFFFFFFC00000000001FFFFFF000000003FFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_27 = 256'hFFFFC000000003FFFFFFFFFFFFFFFFFFFFFE00000000003FFFFFFFFFFFFF07FF;
defparam prom_inst_42.INIT_RAM_28 = 256'hFFE0000000001FFFFFFFFFFFFFC1FFFF3FFFFFFFFFFFFFFFFFF800000000009F;
defparam prom_inst_42.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFF800000000009FFFFF0000000007FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2A = 256'hF4000000001FFFFFFFFFFFFFFFFFFFFFFE000000000FFFFFFFFFFFFFF07FFF8F;
defparam prom_inst_42.INIT_RAM_2B = 256'hF00000000FFFFFFFFFFFFFFC1FFFE3FFFFFFFFFFFFFFFFFFF000000000001FFF;
defparam prom_inst_42.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFF000000000001FFFE0000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2D = 256'h000000007FFFFFFFFFFFFFFFFFFFFFFF0000000FFFFFFFFFFFFFFE03FFF1FFFF;
defparam prom_inst_42.INIT_RAM_2E = 256'h00000FFFFFFFFFFFFFFF81FFFC7FFFFFFFFFFFFFFFFFFFE000000000003FFF00;
defparam prom_inst_42.INIT_RAM_2F = 256'hFFFFFFFFFFFFFE000002000003FF80000000000FFFFFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_42.INIT_RAM_30 = 256'h000001FFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFE07FFC1FFFFFFF;
defparam prom_inst_42.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFF01FFF07FFFFFFFFFFFFFFFFFFFFE000000000013FC00000;
defparam prom_inst_42.INIT_RAM_32 = 256'hFFFFFFFFFFFC0000000000078000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_33 = 256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFC1FFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_34 = 256'hFFFFFFFFFFFFFE03FFF07FFFFFFFFFFFFFFFFFFFFFC000004000007000000000;
defparam prom_inst_42.INIT_RAM_35 = 256'hFFFFFFFFFC000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_36 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FFF81FFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_37 = 256'hFFFFFFFFFFE0FFFE07FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000;
defparam prom_inst_42.INIT_RAM_38 = 256'hFFFFFFFC00000800000000000000010FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFF83FFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3A = 256'hFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFC00000400000000000000041FF;
defparam prom_inst_42.INIT_RAM_3B = 256'hFFFFFC00000400000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3D = 256'hFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFC0000040000000000000000FFFFF;
defparam prom_inst_42.INIT_RAM_3E = 256'hFFFE0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_43 (
    .DO({prom_inst_43_dout_w[29:0],prom_inst_43_dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_43.READ_MODE = 1'b1;
defparam prom_inst_43.BIT_WIDTH = 2;
defparam prom_inst_43.RESET_MODE = "SYNC";
defparam prom_inst_43.INIT_RAM_00 = 256'h555503E9501AAA56C551114D16ABFFFFF9152FFFFFFFAAA7AAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_01 = 256'hAAAA56AAA655403C55AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA555;
defparam prom_inst_43.INIT_RAM_02 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_03 = 256'h5500F9501AAA56805157E45AAFFFFE514FFFFFFFFEAA8AAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_04 = 256'hAAAAAAA955D1156AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9A55555;
defparam prom_inst_43.INIT_RAM_05 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_06 = 256'h40F9502AAA56BC451C816ABFFFE454BFFFFFFFEAA5AAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_07 = 256'hAA9AA554155AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555555;
defparam prom_inst_43.INIT_RAM_08 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_09 = 256'hF9502AAA5AF8504205AAFFFE451FFFFFFFFEAA6AAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_0A = 256'hAA555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555500;
defparam prom_inst_43.INIT_RAM_0B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA6;
defparam prom_inst_43.INIT_RAM_0C = 256'h506AAA96E4041506ABFF944FFFFFFFFFAAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_0D = 256'h5555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555540E9;
defparam prom_inst_43.INIT_RAM_0E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9;
defparam prom_inst_43.INIT_RAM_0F = 256'h6AAA56D084706AAFE543FFFFFFFFFEAEDAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_10 = 256'hAAAAAA9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555540E550;
defparam prom_inst_43.INIT_RAM_11 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAA9AA55;
defparam prom_inst_43.INIT_RAM_12 = 256'hAA56A15381AAA5542FFFFFFFFFAAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_13 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555540E550AA;
defparam prom_inst_43.INIT_RAM_14 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA6AAA;
defparam prom_inst_43.INIT_RAM_15 = 256'h40154D1695542AFFFFFFFFEAA96AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_16 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555540E550AAA9;
defparam prom_inst_43.INIT_RAM_17 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA6AAAAAAAAAAAA9AAAAAA;
defparam prom_inst_43.INIT_RAM_18 = 256'h5570155417EFFFFFFFF0ABB6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_19 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555543E551AAA515;
defparam prom_inst_43.INIT_RAM_1A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAA96AAAAAAAAAAAAAAAA966AAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_1B = 256'h81502BFFAFFFFFFEFAA56AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_1C = 256'hAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555503E541AAAD5856;
defparam prom_inst_43.INIT_RAM_1D = 256'hAAAAAAAAAAAAAAAAAAAA9AA59A6A9AAAAAAAAAAAAAAA9A9AAAAAAAAAA6AAAA9A;
defparam prom_inst_43.INIT_RAM_1E = 256'h9FFFFEBFFFFFF7AAD6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_1F = 256'hAAAAAAAA695AAAAA9AAAAAAAAAAAAAAAAAAAAAAAAAAA555503E552AA36554E00;
defparam prom_inst_43.INIT_RAM_20 = 256'hAAAAAAAAAAAAAAA9AAA5AA99AA95A9A5AAA6AAAAA955AAAAAAAAAA5AA9AAAA6A;
defparam prom_inst_43.INIT_RAM_21 = 256'hFFFBFFFEFEAA95AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_22 = 256'h9A99A5AAAAAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAA5555403A552A9555A92FFFF;
defparam prom_inst_43.INIT_RAM_23 = 256'hAAAAAAAAAAA6AA9955996A66A66669A669696555566A5AA9556A59A559A5AA69;
defparam prom_inst_43.INIT_RAM_24 = 256'hDBFFFFEEB65AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_25 = 256'hA59596AAA96AAAAAAAAAAAAAAAAAAAAAAAAAAAA9555403A546AA5559CCFFFFFF;
defparam prom_inst_43.INIT_RAM_26 = 256'hAAAAAAAAAA555A5555655595565655559555696AAA6A5A5AA565A5A65AA69995;
defparam prom_inst_43.INIT_RAM_27 = 256'hFFEEAA55AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_28 = 256'h555A55569AAAAAAAAAAAAAAAAAAAAAAAAAAAA555540FA55595546C3FFFFFFF7F;
defparam prom_inst_43.INIT_RAM_29 = 256'hAAA696A655555559555565A55595995595595A5595555A556556559556A555A5;
defparam prom_inst_43.INIT_RAM_2A = 256'hEAD96AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_2B = 256'h659555AAAAAAAAAAAAAAAAAAAAAAAAAAAA9955540FA50C15A56FFFFFFFFDEFFF;
defparam prom_inst_43.INIT_RAM_2C = 256'h6555559655555555555555555555A555555555556A65555955A6555565559555;
defparam prom_inst_43.INIT_RAM_2D = 256'h56AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAAAAAAAAAAA9AAAAA;
defparam prom_inst_43.INIT_RAM_2E = 256'h5599565A6AAAAAAAAAAAAAAAAAAAAAAAA555540FA51D10556FFFFFFFE3FFEEB9;
defparam prom_inst_43.INIT_RAM_2F = 256'h5555555955555555556555555556565559555555555556555565655555555555;
defparam prom_inst_43.INIT_RAM_30 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99A5;
defparam prom_inst_43.INIT_RAM_31 = 256'h555A655AAAAAAAAAAAAAAAAAAAAAAAA555503FA523B7556FFFFFF5DFFFAA756A;
defparam prom_inst_43.INIT_RAM_32 = 256'h5555555555555555555555556555559555555555555565555555555555555555;
defparam prom_inst_43.INIT_RAM_33 = 256'hAAAAAAAAAAAAAAAAAAAAAA9AAAAAAA9AAAAAAAAAAAAAAAAAAAAAAAA6A9955555;
defparam prom_inst_43.INIT_RAM_34 = 256'h555AAA6AAAAAAAAAAAAAAAAAAAAA9555503FE8469A55AFFFF6C36FAA9956AAAA;
defparam prom_inst_43.INIT_RAM_35 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_43.INIT_RAM_36 = 256'hAAAAAAAAAAAAAAAAA9AAAAAAAAA9AAAAAAA6AAAAAAAAAA6AAAA6AA5555555555;
defparam prom_inst_43.INIT_RAM_37 = 256'h69A6AAAAAAAAAAAAAAAAAAAAAAA555403FE48F7B56AFEBACF9AAB955AAAAAAAA;
defparam prom_inst_43.INIT_RAM_38 = 256'h5555555555555555555555555555555555555555555555555555555555555559;
defparam prom_inst_43.INIT_RAM_39 = 256'hAAAAAAAAAAAAAAAAA9AAAAAA9AA9AAAA9AAAAA9A9AAA99AA6655555555555555;
defparam prom_inst_43.INIT_RAM_3A = 256'hAAAAAAAAAAAAAAAAAAAAAAAA6555400FE5470C4EA91FFFD6AE455AAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_3B = 256'h555555555555555555555555555555555555555555555555555555555555556A;
defparam prom_inst_43.INIT_RAM_3C = 256'hAAAAAAAAAAA6A55A9AA69AAA999966AA69AA665AA666A5555555555555555555;
defparam prom_inst_43.INIT_RAM_3D = 256'hAAAAAAAAAAAAAAAAAAAAAA5555400FE4C03984A6BFFF7A9155AAAAAAAAAAAAAA;
defparam prom_inst_43.INIT_RAM_3E = 256'h555555555555555555555555555555555555555555555555555555555555556A;
defparam prom_inst_43.INIT_RAM_3F = 256'hAAAAAAAA66956A566595559A9555555555555565555555555555555555555555;

pROM prom_inst_44 (
    .DO({prom_inst_44_dout_w[29:0],prom_inst_44_dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_44.READ_MODE = 1'b1;
defparam prom_inst_44.BIT_WIDTH = 2;
defparam prom_inst_44.RESET_MODE = "SYNC";
defparam prom_inst_44.INIT_RAM_00 = 256'hAAAAA9555555555564000014000000000000155555555555AAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_01 = 256'hAAAAAAAAAAAAA006AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_02 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_03 = 256'hAAAA55555555556400001000000000000155555555556AAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_04 = 256'hAAAAAAAAAA55AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_05 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_06 = 256'hAA5555555555500001400000000000555555555556AAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_07 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_08 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_09 = 256'h555555555550000500000000001555555555556AAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_0A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_0B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_0C = 256'h555555555000140000000001555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_0D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55;
defparam prom_inst_44.INIT_RAM_0E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_0F = 256'h555555500040000000005555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_10 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555;
defparam prom_inst_44.INIT_RAM_11 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_12 = 256'h55554001000000001555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_13 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA555555;
defparam prom_inst_44.INIT_RAM_14 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_15 = 256'h54000400000005555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_16 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555555;
defparam prom_inst_44.INIT_RAM_17 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_18 = 256'h00100000055555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_19 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95555555540;
defparam prom_inst_44.INIT_RAM_1A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_1B = 256'h40000555555555550556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_1C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555555500100;
defparam prom_inst_44.INIT_RAM_1D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_1E = 256'h15555555555554556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_1F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA955555550550500;
defparam prom_inst_44.INIT_RAM_20 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_21 = 256'h5555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_22 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95555555555555555;
defparam prom_inst_44.INIT_RAM_23 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_24 = 256'h5555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_25 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555555555566555555;
defparam prom_inst_44.INIT_RAM_26 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_27 = 256'h5555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_28 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA555555555569555555555;
defparam prom_inst_44.INIT_RAM_29 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_2A = 256'h5556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_2B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55550055555555555555555;
defparam prom_inst_44.INIT_RAM_2C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_2D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_2E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555015555555555555555555;
defparam prom_inst_44.INIT_RAM_2F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_30 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_31 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555444055555555555555555AAA;
defparam prom_inst_44.INIT_RAM_32 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_33 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_34 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA955501005555555429555556AAAAAA;
defparam prom_inst_44.INIT_RAM_35 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_36 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_37 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555440555555416555555AAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_38 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_39 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_3A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55500016554555555556AAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_3B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_3C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_3D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55505117E505555555AAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_3E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_44.INIT_RAM_3F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;

pROM prom_inst_45 (
    .DO({prom_inst_45_dout_w[27:0],prom_inst_45_dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_8),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_45.READ_MODE = 1'b1;
defparam prom_inst_45.BIT_WIDTH = 4;
defparam prom_inst_45.RESET_MODE = "SYNC";
defparam prom_inst_45.INIT_RAM_00 = 256'h235678CB762157777763666799999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_01 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99999999888887766654565;
defparam prom_inst_45.INIT_RAM_02 = 256'h9999999999999999999999999999999999999999999999999999999AAAAAAAAA;
defparam prom_inst_45.INIT_RAM_03 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_04 = 256'h999999A99A99A999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_05 = 256'hAAAAAAAAAAAAA9A9999AA999999999999999999999999999999999999999A999;
defparam prom_inst_45.INIT_RAM_06 = 256'h889886413675746679999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_07 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA999999998888877766554433666;
defparam prom_inst_45.INIT_RAM_08 = 256'h9999999999999999999999999999999999999999999999999AAAAA9AAAAAAAAA;
defparam prom_inst_45.INIT_RAM_09 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_0A = 256'h9A99999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_0B = 256'hAAA9AA999999999999A99999999999999999999999999999999999999999999A;
defparam prom_inst_45.INIT_RAM_0C = 256'h77433456689999999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_0D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA999999999998888777665545666677766;
defparam prom_inst_45.INIT_RAM_0E = 256'h9999999999999999999999999999999999999999999999AAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_0F = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_10 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_11 = 256'h999999999999999AA99999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_12 = 256'h658999999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9A99A9;
defparam prom_inst_45.INIT_RAM_13 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99999999998888777666667777777777865;
defparam prom_inst_45.INIT_RAM_14 = 256'h999999999999999999999999999999999999999A9999AAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_15 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_16 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_17 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_18 = 256'h99A9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9A99A999999;
defparam prom_inst_45.INIT_RAM_19 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAA99999999988888877776666777778888899999;
defparam prom_inst_45.INIT_RAM_1A = 256'h9999999999999999999999999999999999999AAAA9AAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_1B = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_1C = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_1D = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_1E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAAAAAAAAA9999999999999999;
defparam prom_inst_45.INIT_RAM_1F = 256'hAAAAAAAAAAAAAAAAAAAAAA9999999999998888888888888888999999999AAAAA;
defparam prom_inst_45.INIT_RAM_20 = 256'h9999999999999999999999999999999A9A9AAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_21 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_22 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_23 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_24 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAA99999999999999999999999;
defparam prom_inst_45.INIT_RAM_25 = 256'hAAAAAAAAAAAAAAAA9A9A999999999999998888889999999999999AAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_26 = 256'h99999999999999999999999999999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_27 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_28 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_29 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_2A = 256'hAAAAAAAAAAAAAAA9AAAAAAAAAAAAA9AA99999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_2B = 256'hAAAAAAAAAAAAAAAA9999999999999999999999999999AA9AAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_2C = 256'h99999999999999999999999999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_2D = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_2E = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_2F = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_30 = 256'hAAAAAAAAAAAAAAAAAAAAAA9A9999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_31 = 256'hAAAAAAAAAAAA9999999999999999999999999999AAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_32 = 256'h9999999999999999999AAAA9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_45.INIT_RAM_33 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_34 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_35 = 256'h9999999999999999999999999999999999999999999999999999999999999999;
defparam prom_inst_45.INIT_RAM_36 = 256'h0000000000000000000000000000000099999999999999999999999999999999;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_5 (
  .Q(dff_q_5),
  .D(dff_q_4),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_6 (
  .Q(dff_q_6),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_7 (
  .Q(dff_q_7),
  .D(dff_q_6),
  .CLK(clk),
  .CE(oce)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(prom_inst_20_dout[0]),
  .I1(prom_inst_22_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(prom_inst_16_dout[0]),
  .I1(mux_o_12),
  .S0(dff_q_5)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_13),
  .I1(mux_o_14),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(dout[0]),
  .I0(mux_o_16),
  .I1(mux_o_15),
  .S0(dff_q_1)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(prom_inst_20_dout[1]),
  .I1(prom_inst_22_dout[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(prom_inst_4_dout[1]),
  .I1(prom_inst_5_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(prom_inst_6_dout[1]),
  .I1(prom_inst_7_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(prom_inst_17_dout[1]),
  .I1(mux_o_31),
  .S0(dff_q_5)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_3)
);
MUX2 mux_inst_37 (
  .O(dout[1]),
  .I0(mux_o_35),
  .I1(mux_o_34),
  .S0(dff_q_1)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(prom_inst_21_dout[2]),
  .I1(prom_inst_22_dout[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(prom_inst_8_dout[2]),
  .I1(prom_inst_9_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(prom_inst_10_dout[2]),
  .I1(prom_inst_11_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(prom_inst_18_dout[2]),
  .I1(mux_o_50),
  .S0(dff_q_5)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_3)
);
MUX2 mux_inst_56 (
  .O(dout[2]),
  .I0(mux_o_54),
  .I1(mux_o_53),
  .S0(dff_q_1)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(prom_inst_21_dout[3]),
  .I1(prom_inst_22_dout[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(prom_inst_12_dout[3]),
  .I1(prom_inst_13_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(prom_inst_14_dout[3]),
  .I1(prom_inst_15_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(prom_inst_19_dout[3]),
  .I1(mux_o_69),
  .S0(dff_q_5)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_3)
);
MUX2 mux_inst_75 (
  .O(dout[3]),
  .I0(mux_o_73),
  .I1(mux_o_72),
  .S0(dff_q_1)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(prom_inst_43_dout[4]),
  .I1(prom_inst_45_dout[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(prom_inst_23_dout[4]),
  .I1(prom_inst_24_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(prom_inst_25_dout[4]),
  .I1(prom_inst_26_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(prom_inst_39_dout[4]),
  .I1(mux_o_88),
  .S0(dff_q_5)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_89),
  .I1(mux_o_90),
  .S0(dff_q_3)
);
MUX2 mux_inst_94 (
  .O(dout[4]),
  .I0(mux_o_92),
  .I1(mux_o_91),
  .S0(dff_q_1)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(prom_inst_43_dout[5]),
  .I1(prom_inst_45_dout[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(prom_inst_27_dout[5]),
  .I1(prom_inst_28_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(prom_inst_29_dout[5]),
  .I1(prom_inst_30_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(prom_inst_40_dout[5]),
  .I1(mux_o_107),
  .S0(dff_q_5)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_108),
  .I1(mux_o_109),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(dout[5]),
  .I0(mux_o_111),
  .I1(mux_o_110),
  .S0(dff_q_1)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(prom_inst_44_dout[6]),
  .I1(prom_inst_45_dout[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(prom_inst_31_dout[6]),
  .I1(prom_inst_32_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(prom_inst_33_dout[6]),
  .I1(prom_inst_34_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(prom_inst_41_dout[6]),
  .I1(mux_o_126),
  .S0(dff_q_5)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_127),
  .I1(mux_o_128),
  .S0(dff_q_3)
);
MUX2 mux_inst_132 (
  .O(dout[6]),
  .I0(mux_o_130),
  .I1(mux_o_129),
  .S0(dff_q_1)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(prom_inst_44_dout[7]),
  .I1(prom_inst_45_dout[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(prom_inst_35_dout[7]),
  .I1(prom_inst_36_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(prom_inst_37_dout[7]),
  .I1(prom_inst_38_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(prom_inst_42_dout[7]),
  .I1(mux_o_145),
  .S0(dff_q_5)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(dff_q_3)
);
MUX2 mux_inst_151 (
  .O(dout[7]),
  .I0(mux_o_149),
  .I1(mux_o_148),
  .S0(dff_q_1)
);
endmodule //Gowin_pROM4
