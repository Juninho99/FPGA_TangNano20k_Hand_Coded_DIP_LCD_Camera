//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Thu Aug 31 18:51:20 2023

module Gowin_pROM5 (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [15:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire [26:0] promx9_inst_0_dout_w;
wire [8:0] promx9_inst_0_dout;
wire [26:0] promx9_inst_1_dout_w;
wire [8:0] promx9_inst_1_dout;
wire [26:0] promx9_inst_2_dout_w;
wire [8:0] promx9_inst_2_dout;
wire [26:0] promx9_inst_3_dout_w;
wire [8:0] promx9_inst_3_dout;
wire [26:0] promx9_inst_4_dout_w;
wire [8:0] promx9_inst_4_dout;
wire [26:0] promx9_inst_5_dout_w;
wire [8:0] promx9_inst_5_dout;
wire [26:0] promx9_inst_6_dout_w;
wire [8:0] promx9_inst_6_dout;
wire [26:0] promx9_inst_7_dout_w;
wire [8:0] promx9_inst_7_dout;
wire [26:0] promx9_inst_8_dout_w;
wire [8:0] promx9_inst_8_dout;
wire [26:0] promx9_inst_9_dout_w;
wire [8:0] promx9_inst_9_dout;
wire [26:0] promx9_inst_10_dout_w;
wire [8:0] promx9_inst_10_dout;
wire [26:0] promx9_inst_11_dout_w;
wire [8:0] promx9_inst_11_dout;
wire [26:0] promx9_inst_12_dout_w;
wire [8:0] promx9_inst_12_dout;
wire [26:0] promx9_inst_13_dout_w;
wire [8:0] promx9_inst_13_dout;
wire [26:0] promx9_inst_14_dout_w;
wire [8:0] promx9_inst_14_dout;
wire [26:0] promx9_inst_15_dout_w;
wire [8:0] promx9_inst_15_dout;
wire [30:0] prom_inst_16_dout_w;
wire [9:9] prom_inst_16_dout;
wire [30:0] prom_inst_17_dout_w;
wire [9:9] prom_inst_17_dout;
wire [30:0] prom_inst_18_dout_w;
wire [10:10] prom_inst_18_dout;
wire [30:0] prom_inst_19_dout_w;
wire [10:10] prom_inst_19_dout;
wire [30:0] prom_inst_20_dout_w;
wire [11:11] prom_inst_20_dout;
wire [30:0] prom_inst_21_dout_w;
wire [11:11] prom_inst_21_dout;
wire [30:0] prom_inst_22_dout_w;
wire [12:12] prom_inst_22_dout;
wire [30:0] prom_inst_23_dout_w;
wire [12:12] prom_inst_23_dout;
wire [30:0] prom_inst_24_dout_w;
wire [13:13] prom_inst_24_dout;
wire [30:0] prom_inst_25_dout_w;
wire [13:13] prom_inst_25_dout;
wire [30:0] prom_inst_26_dout_w;
wire [14:14] prom_inst_26_dout;
wire [30:0] prom_inst_27_dout_w;
wire [14:14] prom_inst_27_dout;
wire [30:0] prom_inst_28_dout_w;
wire [15:15] prom_inst_28_dout;
wire [30:0] prom_inst_29_dout_w;
wire [15:15] prom_inst_29_dout;
wire [26:0] promx9_inst_30_dout_w;
wire [8:0] promx9_inst_30_dout;
wire [26:0] promx9_inst_31_dout_w;
wire [8:0] promx9_inst_31_dout;
wire [26:0] promx9_inst_32_dout_w;
wire [8:0] promx9_inst_32_dout;
wire [26:0] promx9_inst_33_dout_w;
wire [8:0] promx9_inst_33_dout;
wire [26:0] promx9_inst_34_dout_w;
wire [8:0] promx9_inst_34_dout;
wire [26:0] promx9_inst_35_dout_w;
wire [8:0] promx9_inst_35_dout;
wire [26:0] promx9_inst_36_dout_w;
wire [8:0] promx9_inst_36_dout;
wire [26:0] promx9_inst_37_dout_w;
wire [8:0] promx9_inst_37_dout;
wire [30:0] prom_inst_38_dout_w;
wire [9:9] prom_inst_38_dout;
wire [30:0] prom_inst_39_dout_w;
wire [10:10] prom_inst_39_dout;
wire [30:0] prom_inst_40_dout_w;
wire [11:11] prom_inst_40_dout;
wire [30:0] prom_inst_41_dout_w;
wire [12:12] prom_inst_41_dout;
wire [30:0] prom_inst_42_dout_w;
wire [13:13] prom_inst_42_dout;
wire [30:0] prom_inst_43_dout_w;
wire [14:14] prom_inst_43_dout;
wire [30:0] prom_inst_44_dout_w;
wire [15:15] prom_inst_44_dout;
wire [15:0] prom_inst_45_dout_w;
wire [15:0] prom_inst_45_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire dff_q_7;
wire dff_q_8;
wire dff_q_9;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_49;
wire mux_o_50;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_101;
wire mux_o_102;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_153;
wire mux_o_154;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_205;
wire mux_o_206;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_257;
wire mux_o_258;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_309;
wire mux_o_310;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_361;
wire mux_o_362;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_413;
wire mux_o_414;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_465;
wire mux_o_466;
wire mux_o_484;
wire mux_o_485;
wire mux_o_503;
wire mux_o_504;
wire mux_o_522;
wire mux_o_523;
wire mux_o_541;
wire mux_o_542;
wire mux_o_560;
wire mux_o_561;
wire mux_o_579;
wire mux_o_580;
wire mux_o_598;
wire mux_o_599;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT5 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_0.INIT = 32'h00000001;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(lut_f_0)
);
defparam lut_inst_1.INIT = 4'h8;
LUT5 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_2.INIT = 32'h00000002;
LUT2 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(lut_f_2)
);
defparam lut_inst_3.INIT = 4'h8;
LUT5 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_4.INIT = 32'h00000004;
LUT2 lut_inst_5 (
  .F(lut_f_5),
  .I0(ce),
  .I1(lut_f_4)
);
defparam lut_inst_5.INIT = 4'h8;
LUT5 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_6.INIT = 32'h00000008;
LUT2 lut_inst_7 (
  .F(lut_f_7),
  .I0(ce),
  .I1(lut_f_6)
);
defparam lut_inst_7.INIT = 4'h8;
LUT5 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_8.INIT = 32'h00000010;
LUT2 lut_inst_9 (
  .F(lut_f_9),
  .I0(ce),
  .I1(lut_f_8)
);
defparam lut_inst_9.INIT = 4'h8;
LUT5 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_10.INIT = 32'h00000020;
LUT2 lut_inst_11 (
  .F(lut_f_11),
  .I0(ce),
  .I1(lut_f_10)
);
defparam lut_inst_11.INIT = 4'h8;
LUT5 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_12.INIT = 32'h00000040;
LUT2 lut_inst_13 (
  .F(lut_f_13),
  .I0(ce),
  .I1(lut_f_12)
);
defparam lut_inst_13.INIT = 4'h8;
LUT5 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_14.INIT = 32'h00000080;
LUT2 lut_inst_15 (
  .F(lut_f_15),
  .I0(ce),
  .I1(lut_f_14)
);
defparam lut_inst_15.INIT = 4'h8;
LUT5 lut_inst_16 (
  .F(lut_f_16),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_16.INIT = 32'h00000100;
LUT2 lut_inst_17 (
  .F(lut_f_17),
  .I0(ce),
  .I1(lut_f_16)
);
defparam lut_inst_17.INIT = 4'h8;
LUT5 lut_inst_18 (
  .F(lut_f_18),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_18.INIT = 32'h00000200;
LUT2 lut_inst_19 (
  .F(lut_f_19),
  .I0(ce),
  .I1(lut_f_18)
);
defparam lut_inst_19.INIT = 4'h8;
LUT5 lut_inst_20 (
  .F(lut_f_20),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_20.INIT = 32'h00000400;
LUT2 lut_inst_21 (
  .F(lut_f_21),
  .I0(ce),
  .I1(lut_f_20)
);
defparam lut_inst_21.INIT = 4'h8;
LUT5 lut_inst_22 (
  .F(lut_f_22),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_22.INIT = 32'h00000800;
LUT2 lut_inst_23 (
  .F(lut_f_23),
  .I0(ce),
  .I1(lut_f_22)
);
defparam lut_inst_23.INIT = 4'h8;
LUT5 lut_inst_24 (
  .F(lut_f_24),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_24.INIT = 32'h00001000;
LUT2 lut_inst_25 (
  .F(lut_f_25),
  .I0(ce),
  .I1(lut_f_24)
);
defparam lut_inst_25.INIT = 4'h8;
LUT5 lut_inst_26 (
  .F(lut_f_26),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_26.INIT = 32'h00002000;
LUT2 lut_inst_27 (
  .F(lut_f_27),
  .I0(ce),
  .I1(lut_f_26)
);
defparam lut_inst_27.INIT = 4'h8;
LUT5 lut_inst_28 (
  .F(lut_f_28),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_28.INIT = 32'h00004000;
LUT2 lut_inst_29 (
  .F(lut_f_29),
  .I0(ce),
  .I1(lut_f_28)
);
defparam lut_inst_29.INIT = 4'h8;
LUT5 lut_inst_30 (
  .F(lut_f_30),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_30.INIT = 32'h00008000;
LUT2 lut_inst_31 (
  .F(lut_f_31),
  .I0(ce),
  .I1(lut_f_30)
);
defparam lut_inst_31.INIT = 4'h8;
LUT3 lut_inst_32 (
  .F(lut_f_32),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_32.INIT = 8'h02;
LUT3 lut_inst_33 (
  .F(lut_f_33),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_33.INIT = 8'h08;
LUT5 lut_inst_34 (
  .F(lut_f_34),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_34.INIT = 32'h00010000;
LUT2 lut_inst_35 (
  .F(lut_f_35),
  .I0(ce),
  .I1(lut_f_34)
);
defparam lut_inst_35.INIT = 4'h8;
LUT5 lut_inst_36 (
  .F(lut_f_36),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_36.INIT = 32'h00020000;
LUT2 lut_inst_37 (
  .F(lut_f_37),
  .I0(ce),
  .I1(lut_f_36)
);
defparam lut_inst_37.INIT = 4'h8;
LUT5 lut_inst_38 (
  .F(lut_f_38),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_38.INIT = 32'h00040000;
LUT2 lut_inst_39 (
  .F(lut_f_39),
  .I0(ce),
  .I1(lut_f_38)
);
defparam lut_inst_39.INIT = 4'h8;
LUT5 lut_inst_40 (
  .F(lut_f_40),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_40.INIT = 32'h00080000;
LUT2 lut_inst_41 (
  .F(lut_f_41),
  .I0(ce),
  .I1(lut_f_40)
);
defparam lut_inst_41.INIT = 4'h8;
LUT5 lut_inst_42 (
  .F(lut_f_42),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_42.INIT = 32'h00100000;
LUT2 lut_inst_43 (
  .F(lut_f_43),
  .I0(ce),
  .I1(lut_f_42)
);
defparam lut_inst_43.INIT = 4'h8;
LUT5 lut_inst_44 (
  .F(lut_f_44),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_44.INIT = 32'h00200000;
LUT2 lut_inst_45 (
  .F(lut_f_45),
  .I0(ce),
  .I1(lut_f_44)
);
defparam lut_inst_45.INIT = 4'h8;
LUT5 lut_inst_46 (
  .F(lut_f_46),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_46.INIT = 32'h00400000;
LUT2 lut_inst_47 (
  .F(lut_f_47),
  .I0(ce),
  .I1(lut_f_46)
);
defparam lut_inst_47.INIT = 4'h8;
LUT5 lut_inst_48 (
  .F(lut_f_48),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_48.INIT = 32'h00800000;
LUT2 lut_inst_49 (
  .F(lut_f_49),
  .I0(ce),
  .I1(lut_f_48)
);
defparam lut_inst_49.INIT = 4'h8;
LUT3 lut_inst_50 (
  .F(lut_f_50),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_50.INIT = 8'h20;
LUT6 lut_inst_51 (
  .F(lut_f_51),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14]),
  .I5(ad[15])
);
defparam lut_inst_51.INIT = 64'h0001000000000000;
LUT2 lut_inst_52 (
  .F(lut_f_52),
  .I0(ce),
  .I1(lut_f_51)
);
defparam lut_inst_52.INIT = 4'h8;
pROMX9 promx9_inst_0 (
    .DO({promx9_inst_0_dout_w[26:0],promx9_inst_0_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_0.READ_MODE = 1'b1;
defparam promx9_inst_0.BIT_WIDTH = 9;
defparam promx9_inst_0.RESET_MODE = "SYNC";
defparam promx9_inst_0.INIT_RAM_00 = 288'hEBF5FEFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD6EBF5BADD6EB75B6DB6DB65A26EA;
defparam promx9_inst_0.INIT_RAM_01 = 288'h0C7DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAFF7FBFDFEFF7EBF5FEFD7FBF5FEFD7;
defparam promx9_inst_0.INIT_RAM_02 = 288'hFBFDFEFF7FBFDFEFF7FBFDC31F7FBFDC31F7FBFDFEFF7FBFDFEE18FBFDC31F7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_03 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC31F7FBFDFEFF70C063EFF7FBFDC31F7;
defparam promx9_inst_0.INIT_RAM_04 = 288'h0C063EFF7FB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_05 = 288'h0B85FEE17FB85C6E170B85C2E180C05C2E180C06030170B85C30170C0602E180C0603018;
defparam promx9_inst_0.INIT_RAM_06 = 288'hEBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70BFDC2E17FB85C2E170B85C2E170B85FEE17;
defparam promx9_inst_0.INIT_RAM_07 = 288'hEB75BAFD6EB75B6DD6DB75FADD6EB75BAFD6EB75FAFD7EB75FAFD7EBF5FAFF7EBF5FEFF7;
defparam promx9_inst_0.INIT_RAM_08 = 288'hDB6DB2A2FCB6DB6DB6DB6DB6DB6DB6DBADB6DB6DBADB6DB75B6DB6EB75BADD6EB75B6DD6;
defparam promx9_inst_0.INIT_RAM_09 = 288'hFBF5FEFD7FBF5FEFF7EBF5BAFD7EB75FAFD6EBF5FAFD7EBF5FAFD7EB75FADD7EB6DB6DB6;
defparam promx9_inst_0.INIT_RAM_0A = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5FEFF7FBFDFAFF7;
defparam promx9_inst_0.INIT_RAM_0B = 288'hFBFDFEFF7FBFDFEFF7FBFDC31F7FBFDFEFF7FB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_0C = 288'hFBFDFEFF7FB863EE18FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC31F7;
defparam promx9_inst_0.INIT_RAM_0D = 288'h0C06031F7FB86030180C7DFEE180C7DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_0E = 288'h0B85C2E170B85C3017FB7582FF70B85C30180C06030180C06030180B86030170B85C2E18;
defparam promx9_inst_0.INIT_RAM_0F = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70B85FEFF70B85C2E170B85C2E170B85C2E17;
defparam promx9_inst_0.INIT_RAM_10 = 288'hEB75FADD6EB6DBADD6EB75BADD6EB75BADD6EBF5FAFD7EB75FAFD7EBF5FAFD7FBF5FAFF7;
defparam promx9_inst_0.INIT_RAM_11 = 288'hEB6DBADB6DB6DB6D95DB6DB6DB6DB6DB6DB6DB6DBADB6EB75BADD6EB75BADD7EB75FADD7;
defparam promx9_inst_0.INIT_RAM_12 = 288'hFBFDFEFF7FBFDFEFF7FBF5FEFD7EBFDFEFF7EBFDFAFF7EBF5FAFD7EB75FAFD7FBF5BADD6;
defparam promx9_inst_0.INIT_RAM_13 = 288'hFBFDC31F7FB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FEFF7;
defparam promx9_inst_0.INIT_RAM_14 = 288'h0C7DFEE180C06030180C7DC3018FB863EE180C06030180C063EFF7FBFDC31F7FBFDFEE18;
defparam promx9_inst_0.INIT_RAM_15 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC3018FBFDC30180C7DC3018;
defparam promx9_inst_0.INIT_RAM_16 = 288'h0C05C2E170B85C2E170B86031F7FB86031F70C7DC31F7FBFDFEFF7FB85FEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_17 = 288'h0B85C2E170B85C2E170B85FEE0EE26900D530C06030180C06030180C05C2E170C0603018;
defparam promx9_inst_0.INIT_RAM_18 = 288'hEBF5FEFD7FBFDFEFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE170B85C2E17FB85C2E17;
defparam promx9_inst_0.INIT_RAM_19 = 288'hEB75BADD6EB6DBADD6EB75BADD6EB75BADD6EB75BADD7EBF5BADD7EBF5BAFD7EBF5FEFD7;
defparam promx9_inst_0.INIT_RAM_1A = 288'hEB75FAFD6EB6DBADD6DB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6EB75BADD6EB75BADD6;
defparam promx9_inst_0.INIT_RAM_1B = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAFF7FBFDFEFD7FBF5FEFF7EBFDFAFF7FBF5FAFD7;
defparam promx9_inst_0.INIT_RAM_1C = 288'hFB863EE18FB86031F7FB863EE18FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_1D = 288'h0C06031F70C06030180C06030180C063EFF7FB863EE18FB86030180C7DFEE18FBFDC31F7;
defparam promx9_inst_0.INIT_RAM_1E = 288'hFBFDFEE180C7DFEFF7FB86031F7FBFDFEFF7FBFDFEE18FBFDFEFF70C7DFEE180C7DC3018;
defparam promx9_inst_0.INIT_RAM_1F = 288'h0C06030180B85C2E170B85C2E170B86030180C06030180C7DC31F7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_20 = 288'h0B85C30180C05C2E170B85C2E17FBDD00DA3E271389C4F344C2E180B86030180C0603018;
defparam promx9_inst_0.INIT_RAM_21 = 288'hEBF5FEFF7FBFDFAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70B85C2E17;
defparam promx9_inst_0.INIT_RAM_22 = 288'hDB6DBADD7EBF5BADD6EB6DBADD6DB75BADD6EB75BADD7EB75FAFD7EB75FAFD7EBF5FEFD7;
defparam promx9_inst_0.INIT_RAM_23 = 288'hFBF5FAFD7FBF5FAFD6EBF5FADD6DB6DBADB6DB6DB6DB6DB6DB6DB6EB6DBADD6EB75BADD6;
defparam promx9_inst_0.INIT_RAM_24 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBFDFEFF7FBF5FEFF7EBFDFAFF7;
defparam promx9_inst_0.INIT_RAM_25 = 288'h0C7DFEE18FB863EFF70C7DC30180C06031F7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_26 = 288'hFB86030180C06030180C06030180C06030180C0603018FB86030180C06031F70C7DC3018;
defparam promx9_inst_0.INIT_RAM_27 = 288'hFBFDFEE18FBFDC30180C7DC31F70C7DFEFF7FBFDFEE18FBFDC31F7FB86030180C06031F7;
defparam promx9_inst_0.INIT_RAM_28 = 288'h0C06030180C0602E180C06030170B85C2E170B86030180C06030180C7DC31F7FBFDC2E17;
defparam promx9_inst_0.INIT_RAM_29 = 288'h0B8602E170C05C2E170B85C2E170B85C2FF76570F89A4D1E9349A4E1E938AF20B8603017;
defparam promx9_inst_0.INIT_RAM_2A = 288'hEBF5FEFD7FBF5FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17FB85FEFF70B85C2E17;
defparam promx9_inst_0.INIT_RAM_2B = 288'hEBF5BADB6EB75BAFD6EB75BADD6EB75FADD6EB75BAFD6EBF5BAFD7EB75BAFD7EBF5FEFF7;
defparam promx9_inst_0.INIT_RAM_2C = 288'hFBFDFAFF7FBF5FEFD7FBF5FAFD7EB75FADD6EB75B6DB6DB75B6DB6DB6DBADB6EB75BADD7;
defparam promx9_inst_0.INIT_RAM_2D = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_2E = 288'h0C7DC3018FBFDC31F70C063EE180C0603018FBFDC30180C7DC31F7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_2F = 288'h0C06030180C063EE180C06030180C063EE180C06031F70C06030180C06030180C063EE18;
defparam promx9_inst_0.INIT_RAM_30 = 288'hFBFDC2E170BFDFEFF7FBFDFEFF70C06030180C06031F7FBFDC31F70C06031F70C0603018;
defparam promx9_inst_0.INIT_RAM_31 = 288'h656546E170C0606E180C06030180C06030180C05C2E170B85C2E170B85FEFF70C05C2E17;
defparam promx9_inst_0.INIT_RAM_32 = 288'h0B85FEE170B85C2E170B85C2E170B85C2E170B85C9FC5D268F49A4D271389A4D271349E4;
defparam promx9_inst_0.INIT_RAM_33 = 288'hEBF5BAFD7EBFDFAFD7FBFDFEFD7EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_0.INIT_RAM_34 = 288'hEB75BAFD6EB75BADD6EB75BADD6EB75B6DD6EB75BAFD6EB75BAFD6EBF5BAFD7EBF5FAFD7;
defparam promx9_inst_0.INIT_RAM_35 = 288'hFBFDFEFF7FBFDFEFD7FBF5FAFF7FBF5FAFD7EBF5FADD6EB6DB6DB6DB6DB6DB6DB75B6DD6;
defparam promx9_inst_0.INIT_RAM_36 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FEFF7;
defparam promx9_inst_0.INIT_RAM_37 = 288'h0C0603018FBFDC31F7FB86031F7FB863EE180C063EFF7FB863EE18FBFDFEFF70C7DFEFF7;
defparam promx9_inst_0.INIT_RAM_38 = 288'h0C06030180C06030180C06030180C06030180C063EE180C06030180C06030180C0603018;
defparam promx9_inst_0.INIT_RAM_39 = 288'h0B85C2E170B85C2E170B85FEFF7FB85C2E170BFDC2E170BFDFEE170B85FEE170B85C3018;
defparam promx9_inst_0.INIT_RAM_3A = 288'hD27100A70DADD1A22FDA8602E180C06030180C0602E180C05C2E170B85C2E170B85C2E17;
defparam promx9_inst_0.INIT_RAM_3B = 288'hFB85FEE17FB85C2E170B85C2E170B85C30170B85C2E17FBF59A3E5E270F49C4E269349A4;
defparam promx9_inst_0.INIT_RAM_3C = 288'hEBF5FAFD7EBF5FAFD7EBFDFAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_0.INIT_RAM_3D = 288'hEB75BADB6DB75BADD6EB75BADD6EB75FADD6EB75BAFD7EB6DBADD7EBF5FADD6EB75BAFD6;
defparam promx9_inst_0.INIT_RAM_3E = 288'hFBFDFEFF7FBFDFEFF7FBFDFAFF7EBFDFEFD7EBFDFAFD7EBF5FAFD6EBF5BADB6DB6DB6DB6;
defparam promx9_inst_0.INIT_RAM_3F = 288'hFBFDFEE180C7DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;

pROMX9 promx9_inst_1 (
    .DO({promx9_inst_1_dout_w[26:0],promx9_inst_1_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_1.READ_MODE = 1'b1;
defparam promx9_inst_1.BIT_WIDTH = 9;
defparam promx9_inst_1.RESET_MODE = "SYNC";
defparam promx9_inst_1.INIT_RAM_00 = 288'h0C06030180C06030180C063EE180C063EFF7FBFDC30180C7DFEE180C06031F7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_01 = 288'hFBFDFEE170B85C2E170C06030180C06030180C06030180C06030180C06030180C0603018;
defparam promx9_inst_1.INIT_RAM_02 = 288'h0B85C2FF70BFDC2FF70B85FEFF7FBFDFEFF7FBFDC2E17FB85C2E170BFDC2E170B85C2E17;
defparam promx9_inst_1.INIT_RAM_03 = 288'hD269389A3E1C2B6B9599AA349C4E25B7EC180B85C30170C06030170B85C2E170B85C2E17;
defparam promx9_inst_1.INIT_RAM_04 = 288'hFBFDFEFF70B85FEE17FB85C2E170B85C2E170B85C2FF7FC063AFEE4854FEDF68881789C4;
defparam promx9_inst_1.INIT_RAM_05 = 288'hEBF5FAFD7EBF5FAFD7EBF5FAFD7EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_06 = 288'hDB6DB6DB6EB6DBADD6EB75FADD6EB75BADD7EBF5BADD6EB75FADD6EB75BADD6EB75BAFD7;
defparam promx9_inst_1.INIT_RAM_07 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FEFF7EBF5FEFD7EBFDFEFD7EBFDFADD7EB75BAFB6;
defparam promx9_inst_1.INIT_RAM_08 = 288'h0C7DFEE180C7DC31F7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_09 = 288'h0C06030180C06030180C06030180C06031F70C0603018FB863EFF7FBFDFEFF70C063EFF7;
defparam promx9_inst_1.INIT_RAM_0A = 288'h0B85C2E170BFDC2E170B85C2E170C06030180C06030180C06030180C06030180C0603018;
defparam promx9_inst_1.INIT_RAM_0B = 288'hFBFDC2E170B85C2E170BFDC2FF7FBFDC2FF7FBFDFEFF7FBFDC2E170BFDFEE17FB85C2FF7;
defparam promx9_inst_1.INIT_RAM_0C = 288'hEB0562605E1F0F8626A9ED6A8B0E2E8F87A3D270F8B6CFB7E02E170B85C2E170B85C2E17;
defparam promx9_inst_1.INIT_RAM_0D = 288'hFBFDFEFF7FBFDFEFF70BFDC2E170B85C2E170B85C2E170B85C2E180BB4B89C3E1F14DF34;
defparam promx9_inst_1.INIT_RAM_0E = 288'hEB75BADD6EBF5BAFD6EBF5FAFD7EBF5FAFD7EBF5FAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_0F = 288'hEBF5FADD7EB6DBADD6EB75BADD6EB75BADD6EB75FADD6EB75BADD6EBF5BADD6EB75BAFD6;
defparam promx9_inst_1.INIT_RAM_10 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FAFF7FBFDFEFD7FBFDFAFF7FBF5FAFF7;
defparam promx9_inst_1.INIT_RAM_11 = 288'hFB86031F7FB86031F7FB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_12 = 288'h0C06030180C06031F70C06030180C0603018FB86031F70C0603018FBFDC30180C063EFF7;
defparam promx9_inst_1.INIT_RAM_13 = 288'h0B85C2E170B85C2E170B85C2E170B85C2E170C06030180C7DC30180C06031F70C0603018;
defparam promx9_inst_1.INIT_RAM_14 = 288'h0B85C2E170BFDC2FF7FB85C2E170BFDC2FF70B85FEFF7FBFDFEFF7FBFDFEE17FB85C2FF7;
defparam promx9_inst_1.INIT_RAM_15 = 288'hD268F47C507553ADD599AA3DBD5CA4C84DC4D1E9347C4E1E8F47A3F2B27ADF80C05C2E17;
defparam promx9_inst_1.INIT_RAM_16 = 288'hFBFDFEFF7FBFDFEFF7FBFDC2FF7FB85C2E170B85C2E170B85C2FF81BFDFEFF623F1389A4;
defparam promx9_inst_1.INIT_RAM_17 = 288'hEB75BAFD7EBF5FADD7EBF5FAFD6EBF5FEFD7EBF5FEFF7EBF5FAFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_18 = 288'hFBFDFAFF7EBF5FAFD7EB75BADB6EB75BADB6EBF5BADD7EB75BADB6EB75BAFD6EBF5FADD6;
defparam promx9_inst_1.INIT_RAM_19 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_1A = 288'h0C7DC31F7FB86031F7FBFDFEFF7FB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_1B = 288'h0C06030180C06030180C06030180C06030180C06030180C06030180C06031F70C7DC31F7;
defparam promx9_inst_1.INIT_RAM_1C = 288'hFBFDC2FF7FBFDC2FF70B85C2E170C05C2E170B85C2E170C06030180C063EE180C0603018;
defparam promx9_inst_1.INIT_RAM_1D = 288'hEBFE3EFF7FBFDFEFF70BFDC2FF7FB85C2FF7FBFDFEFF70B85FEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_1.INIT_RAM_1E = 288'hD1E9347A4D268F49A3D1F135973DAFDF2B9417F9389A3D269349A4D268F49C4D1F10CFF6;
defparam promx9_inst_1.INIT_RAM_1F = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FB85C2FF70B85C2E170B85C2E17FB85FDDA4;
defparam promx9_inst_1.INIT_RAM_20 = 288'hEB75FADD6EB75BADD6EBF5FADD7EBF5FAFD7EBF5FAFD7EBFDFAFD7EBF5FAFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_21 = 288'hFBF5FEFF7FBFDFEFF7FBF5FAFD7DB75BADD6EB75BADD6EB75BADD7EB75BADD6EB75BAFD6;
defparam promx9_inst_1.INIT_RAM_22 = 288'hFBFDFEFF7FBFDFEE17FBFDFEFF7FBFDFEFF7FBFDFEFF7EBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_23 = 288'h0C06030180C063EFF7FB86031F70C063EFF7FB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_24 = 288'h0C7DC30180C06030180C06030180C063EE180C06030180C06030180C06030180C0603018;
defparam promx9_inst_1.INIT_RAM_25 = 288'hFB85FEFF7FBFDFEFF7FBFDFEE170B85C2E170C05C2E170B85C2E170C06030180C7DFEE18;
defparam promx9_inst_1.INIT_RAM_26 = 288'hE26B36D753801719D7FBFDFEFF7FBFDFEFF7FBFDFEE17FBFDFEFF7FB85FEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_27 = 288'hBAF9BC7A4E269389A3D269349C3E271111B5EB24121D6BA01B89A3E1E9389C4D271349C3;
defparam promx9_inst_1.INIT_RAM_28 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2FF7FBFDFEE170B85C2E170B85C2FF7;
defparam promx9_inst_1.INIT_RAM_29 = 288'hEB75BAFD7EB75BADD6EB75BAFD6EB75FAFD7EB75FAFD7EBF5FAFD7EBFDFAFF7FBFDFEFD7;
defparam promx9_inst_1.INIT_RAM_2A = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAFD7DB75BADD6EB75BADD6EB75BADD6EB75FADD7;
defparam promx9_inst_1.INIT_RAM_2B = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_2C = 288'h0C06030180C0603018FB86030180C0603018FBFDFEFF7FBFDFEFF7FBFDC31F7FBFDC3018;
defparam promx9_inst_1.INIT_RAM_2D = 288'h0C063EE180C0603018FBFDC3018FBFDC30180C7DFEE180C06030180C063EE180C0603018;
defparam promx9_inst_1.INIT_RAM_2E = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE170B85C2E170B85C30170B85C2E170B85C3018;
defparam promx9_inst_1.INIT_RAM_2F = 288'hD268F8806CA5DAA688E271389A4D675FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_30 = 288'h0B85FEFB6A9A1F49A4D269349A4D271389C4E252B6DD6A9BC89F13EAFDA6845D1E8F89A4;
defparam promx9_inst_1.INIT_RAM_31 = 288'hFBF5FEFF7FBF5FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2FF70BFDC2FF70B85C2E17;
defparam promx9_inst_1.INIT_RAM_32 = 288'hEBF5BADD6EB75FADD6EBF5BAFD7EB75FAFD6EBF5FAFD7EBF5FADD7EBF5FAFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_33 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFD7FBFDFEFF7FBFDFEFD7EB75BADD6EB75BADD6EB75BADD6;
defparam promx9_inst_1.INIT_RAM_34 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70BFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_35 = 288'h0C06030180C06030180C0603018FBFDFEFF7FB86031F7FBFDFEFF7FBFDC31F7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_36 = 288'h0B85C30180C7DC30180C06030180C06031F70C06030180C06030180C063EE180C0603018;
defparam promx9_inst_1.INIT_RAM_37 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70BFDFEE170B85C2E170BFDC2E170B85C2E17;
defparam promx9_inst_1.INIT_RAM_38 = 288'h9981787C3E27139BD5BABC38BC3E1E9349A4E1F101DB6FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_39 = 288'h0B85C2FF7FBAC71B12DB75AA668E269349A4E26938826A9F5B2B1233813C7C3D6DCF6BF7;
defparam promx9_inst_1.INIT_RAM_3A = 288'hEBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70B85FEFF7;
defparam promx9_inst_1.INIT_RAM_3B = 288'hEB75BADD6EB75BADD6EB75BAFD6EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_1.INIT_RAM_3C = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAFF7FBFDFEFF7EBFDFEFF7EB75BADD6EB75BADD6;
defparam promx9_inst_1.INIT_RAM_3D = 288'hFB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_3E = 288'h0C06030180C06030180C06030180C0603018FB863EFF70C06031F7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_1.INIT_RAM_3F = 288'h0B85C2E170B85C2E170B85C2E170B85C2E180C06030180C063EE180C06031F70C0603018;

pROMX9 promx9_inst_2 (
    .DO({promx9_inst_2_dout_w[26:0],promx9_inst_2_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_2.READ_MODE = 1'b1;
defparam promx9_inst_2.BIT_WIDTH = 9;
defparam promx9_inst_2.RESET_MODE = "SYNC";
defparam promx9_inst_2.INIT_RAM_00 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FB85C2E170B85C2E170B85C2E17;
defparam promx9_inst_2.INIT_RAM_01 = 288'hD1F939D73DB7DAA89064DD3AD5364E9389C4E1F1387A3D1E8F49C4F77582FF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_02 = 288'hFBFDC2FF7FBFDFF1B60371389A4D6CD36DD7BA11F49A3D1F1319D6DB4CF59E3E271389C4;
defparam promx9_inst_2.INIT_RAM_03 = 288'hEBF5FAFD7EBFDFEFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2E17;
defparam promx9_inst_2.INIT_RAM_04 = 288'hEBF5BADD7EB75BAFD6EB75BADD6EB75FAFD6EBF5FADD6EB75FAFD7EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_2.INIT_RAM_05 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFD7EB75BADD6;
defparam promx9_inst_2.INIT_RAM_06 = 288'h0C063EFF7FBFDFEFF7FB863EFF7FBFDFEFF7FBFDFEFF7FBF5FEE18FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_07 = 288'h0C0603018FB8603018FB86030180C06030180C06030180C063EE180C7DFEE18FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_08 = 288'h0B85C2E170B85C2E170B85C2FF7FBFDFEFF7EB5D6ABB6FBFDC30180C7DC30180C0603018;
defparam promx9_inst_2.INIT_RAM_09 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70B85C2E170B85C2E17;
defparam promx9_inst_2.INIT_RAM_0A = 288'hE271347A4E1F0F87C5A5DD36DF6FBE566626E1F1387C4E1F1389C3E268F89A4F244B2C17;
defparam promx9_inst_2.INIT_RAM_0B = 288'hFBFDFEFF7FBFDFEFF7FB85BDDC4D1E9349A4E1F105F94CB75EA6E943DCF6DB58881747A4;
defparam promx9_inst_2.INIT_RAM_0C = 288'hFBF5FAFD7EBF5FAFD7EBF5FAFF7FBF5FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_0D = 288'hEB75BADD7EB75BAFD6EB75BAFB6EBF5BADD6EBF5BADD6EB75FADD6EB75FAFD7EB75FAFD7;
defparam promx9_inst_2.INIT_RAM_0E = 288'h0BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_0F = 288'h0C7DFEFF70C7DFEFF7FB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_10 = 288'h0C06030180C06030180C06030180C06030180C06030180C06030180C063EFF7FBFDC31F7;
defparam promx9_inst_2.INIT_RAM_11 = 288'h0B85C30170B85C30170B85C2E17FB85FEFF7EBDD7DEAA44A2514AA967DFF1F8FB8603018;
defparam promx9_inst_2.INIT_RAM_12 = 288'hDAED62595FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2E170B85C2E17;
defparam promx9_inst_2.INIT_RAM_13 = 288'hD278F87C4E1F1389C4E269389C4E2123AB548954F6CB002F8F49C4E271389C3D270F86A8;
defparam promx9_inst_2.INIT_RAM_14 = 288'hFBFDFEFF7FBFDC2FF70BFDFF1F7CAF1749A4D269349A3D269389C4075536DD7DB656656A;
defparam promx9_inst_2.INIT_RAM_15 = 288'hFBF5BAFD7EBF5BAFD7EBF5FAFD7EBF5FAFF7EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_16 = 288'hFBFDFEFF7EBF5BADD7DB75FAFD6EB75BADD6EB75FADD6EB75FADD6EB75BADD6EBF5FADD6;
defparam promx9_inst_2.INIT_RAM_17 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_18 = 288'hFB863EFF7FBFDFEFF7FBFDFEFF7FB863EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_19 = 288'hFBFDC30180C0603018FB86030180C06030180C063EFF70C06030180C06031F70C0603018;
defparam promx9_inst_2.INIT_RAM_1A = 288'hFB85C2E170B85C30170B85C30170B85C2E17FBF5E696D5512493AE34F9C93A6E3AAB6DF7;
defparam promx9_inst_2.INIT_RAM_1B = 288'hF1F1523F6BA8BDC734FBF5FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_2.INIT_RAM_1C = 288'h99C4B6A05E1F1387C4E271389A4E268F49E4C67D76D1227E5269B60B2C78BC3E271347A4;
defparam promx9_inst_2.INIT_RAM_1D = 288'hFBFDFEFF7FBFDFEFF7FB85FEFF7FB85FAD0AD269349A4D269349A4D269347C4E231FAD33;
defparam promx9_inst_2.INIT_RAM_1E = 288'hEBF5FADD7EB75BAFD7FBFDFAFD7FBF5FAFD7FBF5FAFF7FBFDFEFF7FBF5FEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_1F = 288'hFBFDFEFF7FBFDFEFF7EBF5BADD6EB75BADD6EB75B6DD6EB75FADD6EB75FADD6EB75BADD6;
defparam promx9_inst_2.INIT_RAM_20 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_21 = 288'h0C7DC30180C06031F7FB863EFF7FBFDFEFF70C7DFEFF7FBFDFEFF7FBFDFEFF7FB86031F7;
defparam promx9_inst_2.INIT_RAM_22 = 288'h348215796FBFDC30180C06030180C06030180C06030180C06031F70C06030180C0603018;
defparam promx9_inst_2.INIT_RAM_23 = 288'hFBFDFEE170B85C2E170B85C2E170C0602E170B85FEFD748A2914694579FCE92966B821EF;
defparam promx9_inst_2.INIT_RAM_24 = 288'hF271389E4546576D335538D8735EBFDFEFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_25 = 288'h27ED72932BA3476BF6BA09787E4E271389A3E27104D74EB5D1A3A4E2690CF74AA757AC2E;
defparam promx9_inst_2.INIT_RAM_26 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70BF5B9BC4E268F49A4D269349A4D26934804;
defparam promx9_inst_2.INIT_RAM_27 = 288'hEBF5BADD7EB75FAFD7EBF5FAFD7EBF5FAFD7EBFDFAFD7FBF5FEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_28 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7EB75BADD6EB75BADD7EB75BADD6EB75BADD6EBF5FAFD7;
defparam promx9_inst_2.INIT_RAM_29 = 288'hFBFDFEFF7FBFDC2FF7FBFDFEFF7FBFDC2E17FBFDC2FF7FB85FEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_2A = 288'h0C06030180C06030180C0603018FBFDFEFF7FBFDFEE18FB863EFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_2B = 288'hD745226D2A6E9F0E8BCB75FEE18FB86030180C06030180C06030180C06030180C0603018;
defparam promx9_inst_2.INIT_RAM_2C = 288'hFBFDFEFF7FBFDFEE170B85C2E170B85C2E17FB85C2E170BFDF6DAE34A28D228654B2DB4D;
defparam promx9_inst_2.INIT_RAM_2D = 288'h236CE69F6EB7344C2FEB65562C261B0D8734FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_2E = 288'hE1F9111B4CADD16005E191E66F3DAF536805E1F1389A401DB36DB599CAF89E4E271389C4;
defparam promx9_inst_2.INIT_RAM_2F = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7EBFDFEFF7FBFDFEFF7FBCCF29B474F0F49C4E269347A4;
defparam promx9_inst_2.INIT_RAM_30 = 288'hEB75FAFD7EBF5BADD7EBF5FAFD7EBF5F6DD7EBF5FAFD7EBFDFEFF7FBFDFEFF7FBF5FEFD7;
defparam promx9_inst_2.INIT_RAM_31 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5FADD6EB75BAFD6DB75BADD7EB75BAFD7;
defparam promx9_inst_2.INIT_RAM_32 = 288'hFBFDC2FF7FBFDFEE17FBFDC2FF7FB85FEFF7FB85FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_33 = 288'h0C06030180C06030180C06030180C06030180C7DFEFF70C7DFEFF70C7DFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_34 = 288'h28AC96450966381167A359A48A361B8E8BD70C06030180C06030180C06030180C0603018;
defparam promx9_inst_2.INIT_RAM_35 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEE17FB85C2E170B85C2E180B85C2E17FBFDF2B0C552AA59CF;
defparam promx9_inst_2.INIT_RAM_36 = 288'hE271389A4E1F100DB499F57AFD699C2DC6C361B0DC734EBF5FAFD7EBF5FEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_37 = 288'hE1E8F49C4F2B47AB748942BC9C3E279387E5B944F2BF6BA11BC825BA6DB2933F2F9389A4;
defparam promx9_inst_2.INIT_RAM_38 = 288'hEBFDFAFF7EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17FBFDFEFF70B944E553EAED1D384;
defparam promx9_inst_2.INIT_RAM_39 = 288'hEBF5FAFD6EB75BAFD7EB75FADD7EBF5FAFD7EBF5FAFF7FBFDFAFD7EBF5FAFD7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_3A = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EB75FAFD6EB75FAFD6EBF5FADD6;
defparam promx9_inst_2.INIT_RAM_3B = 288'hFBFDFEFF70BFDC2FF7FBFDFEFF7FBFDFEFF70BFDFEE170BFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_3C = 288'h0C06030180C06030180C06030180C06030180C06030180C7DFEE18FBFDC31F7FBFDFEFF7;
defparam promx9_inst_2.INIT_RAM_3D = 288'h65B2954D28A44C2008B361E08C35128D86A2513094704DB7DC2E180C06030180C0603018;
defparam promx9_inst_2.INIT_RAM_3E = 288'hFBFDFEFF7FBFDFEFF7FBFDFEE17FB85FEE170B85C2E170B85C2E180B85C2E17FBF5F6C92;
defparam promx9_inst_2.INIT_RAM_3F = 288'hE271389C4E271389A3E2713C7C495651E75344B8D86C361B0D8714EB75FAFD7EBF5FAFD7;

pROMX9 promx9_inst_3 (
    .DO({promx9_inst_3_dout_w[26:0],promx9_inst_3_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_3.READ_MODE = 1'b1;
defparam promx9_inst_3.BIT_WIDTH = 9;
defparam promx9_inst_3.RESET_MODE = "SYNC";
defparam promx9_inst_3.INIT_RAM_00 = 288'h4954F2BB44471388A9EA652E8F1F270F87C3E270F87C4F27926733DAF57EDD6DAD5319C4;
defparam promx9_inst_3.INIT_RAM_01 = 288'hEBFDFEFF7EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5C1A0C;
defparam promx9_inst_3.INIT_RAM_02 = 288'hEB75FAFD7EB75FAFD7EBF5FADD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_03 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EB75FAFD7EBF5FADD6;
defparam promx9_inst_3.INIT_RAM_04 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17FBFDFEFF70B85FEFF7FBFDFEE17;
defparam promx9_inst_3.INIT_RAM_05 = 288'h0C06030180C06030180C06030180C06030180C06030180C063EE180C06031F7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_06 = 288'hFBFDFAF96493AD94AA34E1E8D467228946A351A8944A361A8944C3A2F5FEFF70C0603018;
defparam promx9_inst_3.INIT_RAM_07 = 288'hEBF5FAFD7EBF5FAFD7FBF5FEFF7FBFDFEFF7FBFDFEFF7FB85C2E170B85C2FF70C05C2FF7;
defparam promx9_inst_3.INIT_RAM_08 = 288'hDAC2B89E4D271389C4E271389C4E271388EADB6556270E330D86C361B0D86F4EBF5BADD7;
defparam promx9_inst_3.INIT_RAM_09 = 288'hFBFDC59EDF6FAD2552DA6D329D5BAD49D5C4D1F0F87A3E1F0F89A3E26938806DA54F2994;
defparam promx9_inst_3.INIT_RAM_0A = 288'hEBF5FEFD7FBFDFEFF7FBFDFEFF7FBF5FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_0B = 288'hEB75BADD7EB75BADD6EB75FADD6EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFF7FBF5FEFF7;
defparam promx9_inst_3.INIT_RAM_0C = 288'hFBFDC2FF7FBFDFEE17FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5BADD6;
defparam promx9_inst_3.INIT_RAM_0D = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70BFDFEE170BFDC2FF7FB85FEE17;
defparam promx9_inst_3.INIT_RAM_0E = 288'h0C7DC30180C06030180C06030180C06030180C06030180C06030180C063EE180C0603018;
defparam promx9_inst_3.INIT_RAM_0F = 288'h0B8602FF7FBFDFAFD6CB2C9D6AB24D9A488341B0904C25128944A23118906E461F5BEFF7;
defparam promx9_inst_3.INIT_RAM_10 = 288'hDB75BADD6EB75BAFD7EBF5FAFD7EBF5FEFF7FBFDFEFF70BFDFEE170B85C2E170B85C2E17;
defparam promx9_inst_3.INIT_RAM_11 = 288'hEB6D79DADCA75AA846E279389C3E271389A4E279123B69A3AF8C6F1430D86C361B0DC755;
defparam promx9_inst_3.INIT_RAM_12 = 288'hFBFDFEFF7FBFDEADEDE67B019CA59D4FAB74A971787C4E1F0F87C3E270F87A3E2793C929;
defparam promx9_inst_3.INIT_RAM_13 = 288'hFBF5FAFD7FBF5FEFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_14 = 288'hEBF5BADD6EB75BAFD7EB75FADD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5BAFD7FBF5FAFF7;
defparam promx9_inst_3.INIT_RAM_15 = 288'hFBFDFEFF7FBFDC2FF7FB85FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_16 = 288'h0C0603018FB8603018FBFDFEFF7FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEE17FBFDFEE17;
defparam promx9_inst_3.INIT_RAM_17 = 288'hB334FADF7FBFDC30180C06030180C0602E180C06031F7FBFDC30180C06030180C0603018;
defparam promx9_inst_3.INIT_RAM_18 = 288'h0B85C2E170B85FEFF7FBFDFEFD7DB5D5648A92C9544A25128944A35118882E4724164B24;
defparam promx9_inst_3.INIT_RAM_19 = 288'h71C0C1F95DB6DB6DD6EB75BADD6EB75FAFD7EBF5FEFF7FBFDFEFF70BFDC2E170B85C2E17;
defparam promx9_inst_3.INIT_RAM_1A = 288'hF1815E5D7CAC48CF33DA5CF29D7DA01B89C4E271389E33465B6AD371B0F0A4F44B8D86C3;
defparam promx9_inst_3.INIT_RAM_1B = 288'hFBFDFEFF7FBFDFEFF7FBFDFF1ECF67B3D9ECF64B52133EB03BCBE3D1F0F89C3E271387C4;
defparam promx9_inst_3.INIT_RAM_1C = 288'hEBF5FAFF7FBFDFAFD7FBF5FEFD7FBFDFEFF7FBFDFEFF7FBF5FEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_1D = 288'hFBFDFEFF7EB75FADD7EB75BAFD6EBF5FAFD7EB75FAFD7EB75BAFD7EB75FADD7EB75FAFF7;
defparam promx9_inst_3.INIT_RAM_1E = 288'hFBFDFEE17FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_1F = 288'h0C7DC30180C06030180C06030180C7DC2E17FBFDFEFF7FBFDFEFF70BFDC2FF7FBFDFEE17;
defparam promx9_inst_3.INIT_RAM_20 = 288'h524964B46B359C21D6FBFDC30180C06030180C0602E180C0603018FBFDFEFF70C7DC3018;
defparam promx9_inst_3.INIT_RAM_21 = 288'h0B85C2E170B85C2E170B85C2E17FBFDFEFF7EBEDAEA9255C0D44825128D4461314164A81;
defparam promx9_inst_3.INIT_RAM_22 = 288'h75B0D86C3C30BDA4B2DB6DB6DB6DB6DB6DD6EB75BAFD7EBF5FEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_3.INIT_RAM_23 = 288'hE1F0F89E484EDB6D53D6713C7E4E18166553BA05F2A47F2713C9CDEBD535CC25130E086F;
defparam promx9_inst_3.INIT_RAM_24 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEF2FF6FB3D9ECF67ADA090AA6DBEC4FF270F87C3;
defparam promx9_inst_3.INIT_RAM_25 = 288'hEBFDFAFD7FBF5FAFD7FBF5FEFF7FBFDFAFF7FBFDFEFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_26 = 288'hFBFDFEFF7FBFDFEFF7EBF5BADD6EBF5BADD6EB6DBADD7EBF5BAFD6EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_3.INIT_RAM_27 = 288'hFBFDFEFF7FBFDFEFF7FBFDC2E17FBFDFEFF7FBFDC2FF70B85FEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_28 = 288'h0B85FEE170B85FEE170B85FEFF7FB86030180C05FEE17FB85FEFF7FBFDC2FF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_29 = 288'h92A09C946A3496CC8292B8ECD2DEBFDFEFF70C06030180C06030170B85FEFF7FB85C2E17;
defparam promx9_inst_3.INIT_RAM_2A = 288'hFBFDFEFF7FB85C2E170B85C2E170B85C2E170BFDFEFF7FBF5F6D5549699C6A261209CB05;
defparam promx9_inst_3.INIT_RAM_2B = 288'h5130E062FA630DC72C487B9876DCB6DB6DB6DB6DB6DD6EB75BADD6EB75FEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_2C = 288'hEB0BFC9C4F27100AB1DB6D665C60271389C4E271389E6A95D2EBD6CADB2A79579D9544A3;
defparam promx9_inst_3.INIT_RAM_2D = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFB7067B7D9ECF67B1224FE5D3AA7D6;
defparam promx9_inst_3.INIT_RAM_2E = 288'hEBF5FAFF7EBF5FAFD7EBF5FAFF7EBFDFAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_2F = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7EB75BADD7EBF5FADD6EBF5FAFD6EB75FAFD7EB75FAFD7;
defparam promx9_inst_3.INIT_RAM_30 = 288'hFBFDC2FF7FB85FEFF7FBFDFEE17FBFDFEFF7FBFDC2FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_31 = 288'hFB85C2FF70B85C2E170B85C2E170B85C31F70C0603018FBFDFEFF7FBFDC2E17FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_32 = 288'h20B928B6641D1A4D25A29868D66A35168D4524EDBEFF70C06030180C06030170B85C2E18;
defparam promx9_inst_3.INIT_RAM_33 = 288'hFBFDFEE17FBFDC2FF7FBFDC2E170B85C2E170B85FEFF7FBFDFEFF7FBF5F6D959A03ECAE3;
defparam promx9_inst_3.INIT_RAM_34 = 288'h5130D46A36130E062F2840C1EB11438DC90CCB65B2D96DB6DB6DB6DB75BADD6EBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_35 = 288'h15FB7D7B0BA757AFCC02B236BB5AA0BFC9C3E270F89E4E271389C3E27962394BA7DF6A91;
defparam promx9_inst_3.INIT_RAM_36 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF78AFAFD9EDF67B1586E;
defparam promx9_inst_3.INIT_RAM_37 = 288'hEB75FAFD7EBF5BAFD7EBFDFAFD7EBF5FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_3.INIT_RAM_38 = 288'h0BFDC2FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5BADD6EB75BADD6EB75BADD7EBF5BAFD7;
defparam promx9_inst_3.INIT_RAM_39 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEE17FBFDFEFF70BFDFEFF7FBFDC2E17FBFDFEFF7FBFDC2FF7;
defparam promx9_inst_3.INIT_RAM_3A = 288'h0B8602E170B85C2E170C05C2E170B85C2E170B85C30180C06030180C05FEE17FBFDC2FF7;
defparam promx9_inst_3.INIT_RAM_3B = 288'hBABCC21454120A8D66B351A8CE4B35148482A34128D66B37232BF7FBFDC2E170B8602E17;
defparam promx9_inst_3.INIT_RAM_3C = 288'hEBFDFEFF7FBFDFEFF7FBFDFEFF7FB85C2FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FAFB6;
defparam promx9_inst_3.INIT_RAM_3D = 288'hCA941E6E361B0D86C361B0DC60F480BCE0C371B0D86EBBAE572B96CB65B6DB6DB75BADD7;
defparam promx9_inst_3.INIT_RAM_3E = 288'hF6F33D690D77B7D9EDF67C729B6EB75B6B333370F87C4E270F89C4E1F13C9C4E27100B75;
defparam promx9_inst_3.INIT_RAM_3F = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFD6EB347E1EC;

pROMX9 promx9_inst_4 (
    .DO({promx9_inst_4_dout_w[26:0],promx9_inst_4_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_9),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_4.READ_MODE = 1'b1;
defparam promx9_inst_4.BIT_WIDTH = 9;
defparam promx9_inst_4.RESET_MODE = "SYNC";
defparam promx9_inst_4.INIT_RAM_00 = 288'hEBF5BAFD6EBF5FAFD7EBF5FAFD7EBF5FEFD7EBF5FAFD7EBFDFEFF7FBF5FEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_01 = 288'h0BFDC2FF7FBFDC2FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EB75BADD7EBF5FAFD7EB75FADD6;
defparam promx9_inst_4.INIT_RAM_02 = 288'hFB85FEFF70BFDFEFF7FBFDFEFF7FB85C2FF7FB85C2FF7FB85C2E17FB85FEFF7FBFDFEE17;
defparam promx9_inst_4.INIT_RAM_03 = 288'h0B8602E170B85C31F70B85C30180B85C30170B85C2E170B86030180C0603018FB85C2FF7;
defparam promx9_inst_4.INIT_RAM_04 = 288'hFBFDFAFD6DB65668D3185B7CF86A359A8D46929068D4692D9A08A3A2D174F96FB85C2E17;
defparam promx9_inst_4.INIT_RAM_05 = 288'hDB75BADD6EB75FEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_06 = 288'hE221F6B74588BD21A661A8986C361B0E074C688BD86C361B0D868ABADD72B75CB65B6DB6;
defparam promx9_inst_4.INIT_RAM_07 = 288'hFB82C62D1C7FB3985007733980DE6FB3D892BA5D3684FE278F89C4E1F0F87C3E270F89E3;
defparam promx9_inst_4.INIT_RAM_08 = 288'hEBF5FEFF7FBF5FEFF7FBFDFAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5BEFF6;
defparam promx9_inst_4.INIT_RAM_09 = 288'hEB75BAFD7EBF5FAFD6EB75FADF7EBF5FAFD7FBF5FAFD7EBFDFAFD7EBF5FEFF7FBF5FEFF7;
defparam promx9_inst_4.INIT_RAM_0A = 288'hFBFDFEE17FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EB75FAFD7EBF5FAFD7;
defparam promx9_inst_4.INIT_RAM_0B = 288'hFB85C2E170B85FEFF70BFDFEFF7FBFDFEFF7FB85FEFF7FB85FEFF7FB85FEFF7FB85FEFF7;
defparam promx9_inst_4.INIT_RAM_0C = 288'hAAFDFEE17FB85C2E170B86030170C05C30180B85C30170B85C2E170B85C30180C0603018;
defparam promx9_inst_4.INIT_RAM_0D = 288'hFBFDFEFF7FBFDFEFD7FBF5B2D959A2CB5C69C351ACCC3A2D1A8D465198A8D46A351A4B87;
defparam promx9_inst_4.INIT_RAM_0E = 288'hCB65B6DB6DB6DBADD6EB75FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_0F = 288'hE1F1387E406ED666C961739228961B0D44C361B8C1E0E58A89C4C361B0DC628AADD6EB95;
defparam promx9_inst_4.INIT_RAM_10 = 288'hFBF5BEFD7EAD3C1BCB493469C8C2712F9BECE6737DBCC69BCAA994EAD2FC9C3E270F89C4;
defparam promx9_inst_4.INIT_RAM_11 = 288'hFBFDFEFF7EBFDFEFD7FBF5FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_12 = 288'hEB75BAFD6EB75BADD7EBF5BAFF7EB75FAFD7EBF5FAFD7FBF5BEFD7FBF5FAFD7EBF5FEFF7;
defparam promx9_inst_4.INIT_RAM_13 = 288'hFB85C2E170B85C2FF70BFDFEFF70BFDFEFF70BFDFEE17FBFDFEFF7FBFDFEFF7EB75BADD6;
defparam promx9_inst_4.INIT_RAM_14 = 288'h0C06030170B85C2E170B85FEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17FBFDFEE170BFDFEFF7;
defparam promx9_inst_4.INIT_RAM_15 = 288'h82C128D46C3BCFEFF7FB85C2E170B85C2E180B85C2E180B85C2E170B85C2E170B85C3017;
defparam promx9_inst_4.INIT_RAM_16 = 288'hDB556CB048675BAFD7EBFDFEFF7FBF5F6DB6CAD51E7EF5561ACD46B35164B25A2D98C4E4;
defparam promx9_inst_4.INIT_RAM_17 = 288'hAAD56EB75CAE572DB6DB75BADD6EBF5FAFD7FBFDFEFF7FBFDFEFF7FBFDFAFD6EB5D52375;
defparam promx9_inst_4.INIT_RAM_18 = 288'hE279389C4E1F0C8F53DA3CA488261BA8A18D61B0D86C3C294163EEE730DC6E371B8DC669;
defparam promx9_inst_4.INIT_RAM_19 = 288'hFBFDFEFF7FBFDFADD6EB6581BECF672D64F137FBF59CDF67B7DBED66BC8208C99E5769AB;
defparam promx9_inst_4.INIT_RAM_1A = 288'hEBF5FEFD7EBFDFEFF7FBF5FAFF7FBFDFEFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_1B = 288'hEB6DBAFD7EBF5BAFD7EBF5BAFD7EB75FADD7EBF5FAFD7EBF5FAFD6EBF5FAFF7FBF5FAFD7;
defparam promx9_inst_4.INIT_RAM_1C = 288'hFB85FEE170BFDFEE17FB85FEE17FBFDFEE17FBFDFEFF70BFDFEFF7FBFDC2FF70BFDFEFF7;
defparam promx9_inst_4.INIT_RAM_1D = 288'h0B8602E170B85C2E170BFDC2FF7FBFDFEFF7FBFDC2FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_1E = 288'h414968D86B351989465161D65D7FB85C2E170B85C2E170B85C2E170B85C2E180B85C2E17;
defparam promx9_inst_4.INIT_RAM_1F = 288'hC730E08C35530E4986824B2CAE351043ADD7FBFDFAFD6DB65AA8F3082AB0D46A351A8B26;
defparam promx9_inst_4.INIT_RAM_20 = 288'h71B8ECAF2AA552AB75BAE572DB6DB75BADD6EBF5FAFD7EBFDFEFF7FBFDFAFD7EBF5B6D95;
defparam promx9_inst_4.INIT_RAM_21 = 288'hE64BA27B5DADAFCBE4F24AF6B530720986C36181C5E3061B0D86EB488BD440E17B8D86C3;
defparam promx9_inst_4.INIT_RAM_22 = 288'hFBFDFEFF7FBFDFEFF7EB75BEFD6EB758160CF6FB3D82B69A431FCCE67B7DBEDF5BC923EC;
defparam promx9_inst_4.INIT_RAM_23 = 288'hEBF5FEFD7EBFDFAFD7EBF5FAFF7EBFDFEFD7EBFDFEFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_24 = 288'hFBFDFEFF7EB75BAFD7EB75FAFD6EB75BADD7EB75BAFD7EBF5FAFD7EBF5FAFD7EBF5FEFF7;
defparam promx9_inst_4.INIT_RAM_25 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEE170B85FEE170B85FEFF70BFDFEFF7FBFDFEFF7FBFDC2E17;
defparam promx9_inst_4.INIT_RAM_26 = 288'h0B8602E170B85C2E17FB85C2FF7FB85FEFF70B85C2FF7FBFDFEFF7FBFDFEFF7FB85FEFF7;
defparam promx9_inst_4.INIT_RAM_27 = 288'h92D9A8CA3B359A8D2520516CD67B3E1F0E31FBFDFEE170B85C2E170B85C2E180C05C2E17;
defparam promx9_inst_4.INIT_RAM_28 = 288'hBAE19C78661A0A48C33098609046190587A692A8A68CB75EDBAFD7EBEDB6D75798C197A6;
defparam promx9_inst_4.INIT_RAM_29 = 288'h3830D86E371923DC0F9A552AB75BAE576DB6DB75BADD6EBF5FAFD7EBF5FEFD7EBF5FADB6;
defparam promx9_inst_4.INIT_RAM_2A = 288'hF6349A40CE6F37992E996D7282E8965225C55130D86C361C939C7171C105EB19630DC62F;
defparam promx9_inst_4.INIT_RAM_2B = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFD6EB75BADD6EB6D9EBEDE67B399EC5613DA271F5F37D9ED;
defparam promx9_inst_4.INIT_RAM_2C = 288'hEBFDFAFD7EBF5FAFD7EBFDFAFD7FBF5FAFD7FBF5FAFD7EBFDFEFF7EBF5FEFF7FBF5FAFF7;
defparam promx9_inst_4.INIT_RAM_2D = 288'hFBFDC2FF7FBFDFEFF7EB75BADD6EB75BADD7EBF5FADF7EBF5FADD6EBF5FAFD7EBF5FEFD7;
defparam promx9_inst_4.INIT_RAM_2E = 288'hFBFDC2FF7FBFDFEFF7FBFDC2E17FBFDC2E170B85FEFF70B85C2FF70BFDFEFF70BFDFEFF7;
defparam promx9_inst_4.INIT_RAM_2F = 288'h0B85C2E180B85C2E170B85C2E170B85C2E170B85C2E17FBFDFEFF7FB85FEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_30 = 288'hBAC4CA10BD3D16CD66A35990366B3391C98610E1ECD87E7FDFEFF7FB85C2E170B85C3018;
defparam promx9_inst_4.INIT_RAM_31 = 288'hEBF5B6D759238F0D043098504A24128986C36198504827190587048230B6DF7EBEDBADB6;
defparam promx9_inst_4.INIT_RAM_32 = 288'h61B0DC62F38309C703D75B6076D9A4D2A955BAE5B6DB6DB75BADD6EB75FAFD7EBF5FAFD7;
defparam promx9_inst_4.INIT_RAM_33 = 288'h791C799ECF6E41E4ADE6F3799CCE6DBE6795CA34544A351B0D86C361B8F5A91488BD6344;
defparam promx9_inst_4.INIT_RAM_34 = 288'hFBFDFEFF7FBFDFEFF7FBFDFAFF7FBFDFEFD6EB75BADD6EB75B2DEBF673399ECF59C09DAA;
defparam promx9_inst_4.INIT_RAM_35 = 288'hEBF5FAFD7FBFDFAFD7EBF5FAFD7EBF5FEFD7EBF5FEFF7FBFDFEFD7EBF5FAFD7EBFDFAFD7;
defparam promx9_inst_4.INIT_RAM_36 = 288'hFBFDFEFF7FBFDC2E17FBFDFEFF7EB75BADD7EBF5FAFD6EBF5FAFD6EBF5BAFD7EBF5BAFF7;
defparam promx9_inst_4.INIT_RAM_37 = 288'hFB85FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2E17FBFDFEE17FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_38 = 288'h0B85C2E170B8602E170B86030170B85C2E170B85C2E17FBFDC2E170BFDFEFF7FBFDFEFF7;
defparam promx9_inst_4.INIT_RAM_39 = 288'h82023AFB6DB5D626718669E8D86B361ACD6772D9D8786C361A8D87C3D37EFD7FB85C2FF7;
defparam promx9_inst_4.INIT_RAM_3A = 288'hEBCD3ADD6DB655E6AA6198504C34130DC76585B2C0FE744F9DC6E371984C2C3A29874CE4;
defparam promx9_inst_4.INIT_RAM_3B = 288'h588BD86E361B0DC60F3838E884F24412098D8A4D2A975CAE5B6DB6EB75BADD7EBF5FAFD6;
defparam promx9_inst_4.INIT_RAM_3C = 288'hE59445FEA068AE2451E60AE2652F6F339BCCE673797137963586C361B0D86C361B8F1890;
defparam promx9_inst_4.INIT_RAM_3D = 288'hEBFDFEFF7FBF5FAFF7FBFDFEFF7FBFDFAFF7FBFDFEFF7EB75BADD6EB6DB6B75F57B399CC;
defparam promx9_inst_4.INIT_RAM_3E = 288'hEB75FAFF7EBF5FAFF7EBFDFAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFF7EBF5FEFF7;
defparam promx9_inst_4.INIT_RAM_3F = 288'h0BFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEFF7EB75BADD7EB75BAFD6EBF5FADD7EBF5FADD7;

pROMX9 promx9_inst_5 (
    .DO({promx9_inst_5_dout_w[26:0],promx9_inst_5_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_11),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_5.READ_MODE = 1'b1;
defparam promx9_inst_5.BIT_WIDTH = 9;
defparam promx9_inst_5.RESET_MODE = "SYNC";
defparam promx9_inst_5.INIT_RAM_00 = 288'h0B85FEFF7FBFDFEFF7FB85FEFF7FBFDFEE17FBFDC2E170B85C2E17FB85C2FF7FBFDFEE17;
defparam promx9_inst_5.INIT_RAM_01 = 288'hFBFDFEE170B85C2E170B85C2E170B85C2E170B85C30170B85C2E170BFDC2FF7FB85FEFF7;
defparam promx9_inst_5.INIT_RAM_02 = 288'h411054586C3411A5B6DB65AEB1338D33CF66B3E1E4B87C361B0E414161DC966B3E1D97D6;
defparam promx9_inst_5.INIT_RAM_03 = 288'hEB75BADD6EB75B6D96BAAC986E38230D44E3555B75C10492C964923883E588A24F198682;
defparam promx9_inst_5.INIT_RAM_04 = 288'h61E9B9AD185A8986C371B8E09AD381209EE382411C76D8A4D2A995CB6DB6DB6DB75BADD6;
defparam promx9_inst_5.INIT_RAM_05 = 288'h68F3F97ECF622CDFAFE67B3DACCA9FBE24D1F5F3399CCE66B35B6E789C186C361B0D86C3;
defparam promx9_inst_5.INIT_RAM_06 = 288'hFBF5BAFD7EBF5FEFF7EBD56DC10DB7DFEFF7FBFDFAFD7FBF5BEFD6EB75BADD6DB6DB6B74;
defparam promx9_inst_5.INIT_RAM_07 = 288'hEBF5FAFD7EBF5FAFD7EBF5BEFD7EBF5FAFD7EBF5FAFD7EBF5FAFF7EBF5FAFD6EBF5FEFD6;
defparam promx9_inst_5.INIT_RAM_08 = 288'h0BFDFEE17FBFDFEE17FB85FEFF7FBFDC2FF70BFDFEFF7DB75BADD6EB75BADD7EB75BAFD7;
defparam promx9_inst_5.INIT_RAM_09 = 288'hFB85FEFF7FB85C2FF7FBFDFEFF7FBFDFEFF7FBFDFEE17FBFDC2E170B85C2E170B85C2FF7;
defparam promx9_inst_5.INIT_RAM_0A = 288'h82C96CE49DB7DFEFF7FBFDC2E170B85C30170C05C2E170B85C2E170B85C2FF7FBFDC2E17;
defparam promx9_inst_5.INIT_RAM_0B = 288'h38EB851459241104A39298554D2DB6DB6D7589A4699E7B2E1B0F86C3B11C787C3D9B0D05;
defparam promx9_inst_5.INIT_RAM_0C = 288'hDB75BADD6EBF5FADD6DB6DB6D759A0A0C304A2A8BCF0C0834E2954AADD6AB55AACD226D3;
defparam promx9_inst_5.INIT_RAM_0D = 288'h61B0D86C3E38BF5A916130D86E371B8DC72C0713DC6E471C12096D8A552EB96CB6DB6DB6;
defparam promx9_inst_5.INIT_RAM_0E = 288'hDB6DB2BB5F52C9614EE5FA8E250D5FB7D9EDF62CAE64E56F339BCCE6F33980A792C586C3;
defparam promx9_inst_5.INIT_RAM_0F = 288'hEBEDB6D4D257C3AFD6EBF5FEFF766315CAC562827AFD7FBFDFAFF7EB75BEFD6EB75BADB6;
defparam promx9_inst_5.INIT_RAM_10 = 288'hEB75BAFD7EBFDFAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FEFD7EBFDFAFD7EBF5FADD7;
defparam promx9_inst_5.INIT_RAM_11 = 288'hFBFDFEFF70BFDFEE170B85FEFF7FBFDC2FF7FBFDFEFF7FBFDFEFF7EB75BADD6EB75BADD6;
defparam promx9_inst_5.INIT_RAM_12 = 288'h0B85C2FF70B85FEFF7FBFDFEE17FBFDC2FF7FBFDFEFF7FBFDC2FF7FBFDFEFF7FBFDC2FF7;
defparam promx9_inst_5.INIT_RAM_13 = 288'hC3A054786B3D9ACD66F46DBEFF7FBFDFEE170B85C2E170B85C2E170B85C2E170B85C2E17;
defparam promx9_inst_5.INIT_RAM_14 = 288'hDB65AEB75AA44D6430D72AA08C330B8E090471E5BADB6BACD1236D0459B0D873159ECF67;
defparam promx9_inst_5.INIT_RAM_15 = 288'hCB6DB6DB6DB75BADD6EBF5BADB6DB6DAEB5407B8DC882514139EB29A5D72BB6DB6DB6DB6;
defparam promx9_inst_5.INIT_RAM_16 = 288'h88B4584C361B8DC74C287B8609003B0DC6E361C12887037B0A08E371C12096D9A5D72D96;
defparam promx9_inst_5.INIT_RAM_17 = 288'hEB75BADD6DB6D76B9476F3452B157CB8604FF57B3D9CCF68389911B9BCF97CDE673399EB;
defparam promx9_inst_5.INIT_RAM_18 = 288'hEBF5FAFD7EBE5A0CE662A918A72FBFDFAFD7E431548A462397AFF7EBFDF2DC88351A29D6;
defparam promx9_inst_5.INIT_RAM_19 = 288'hEBF5BAFD7EB75BADD6EB75FAFD6EBFDFAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_5.INIT_RAM_1A = 288'hFBFDC2E170B85C2E170BFDFEE170BFDC2E170BFDFEFF7FBFDFEFF7FBFDFEFF7EB75BADD7;
defparam promx9_inst_5.INIT_RAM_1B = 288'h0B85C2E170B85FEFF7FBFDC2E17FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_5.INIT_RAM_1C = 288'hC3E1ACE8282D9ACCE4A328DCB86B361EABD7EBFDFEFF7FBFDFEE170BFDC2E170B85C2E17;
defparam promx9_inst_5.INIT_RAM_1D = 288'hEB75FADD6EB75BADB6DB656AB347994619A68230E4B244165B6DD6DB5D66891C68230D67;
defparam promx9_inst_5.INIT_RAM_1E = 288'hCB65B6DB6DB6DB6DB6DB75BADD6EB75BADB6DB65AA8D3514930EE4925B52534CAEDB6DD6;
defparam promx9_inst_5.INIT_RAM_1F = 288'hE673399AC89347CCC361C90A091E33901E7095B8DC6E3720A0E22F17A89C6E371C130AD2;
defparam promx9_inst_5.INIT_RAM_20 = 288'h72A914AF4EB75BADD6DB6D72D959A72FD9CC05AC561EEE7FB3D9EDF67B7D9127954EA92F;
defparam promx9_inst_5.INIT_RAM_21 = 288'hEBF5FAFD7EBF5FAFD7EBCD1CCC46231589E8EBFDFAFD682A9148A452317ADD6EBF5B90C5;
defparam promx9_inst_5.INIT_RAM_22 = 288'hEB75BADD7EB75BAFD7EB75BAFD6EBF5FAFD7EBF5FAFD7EBFDFAFD7EBF5FAFD7EBF5FAFD6;
defparam promx9_inst_5.INIT_RAM_23 = 288'hFBFDFEFF7FBFDC2FF70BFDFEE17FB85FEFF70B85FEE170B85C2E17FB85C2FF7FBFDFEFF7;
defparam promx9_inst_5.INIT_RAM_24 = 288'hFBFDFEE170B85FEE170B85C2FF7FBFDFEFF7FBFDC2E17FBFDFEFF70B85C2FF7FBFDFEE17;
defparam promx9_inst_5.INIT_RAM_25 = 288'h596381166B359A4B66B34970C839361A8D46B330F4EF3EB6DB6DD7FBFDFEFF7FB85C2E17;
defparam promx9_inst_5.INIT_RAM_26 = 288'hCB75B6DD6EBF5FAFD7EBF5FAFD7EB6DB6D96BACD1658DB2B0CC24130C118775DB6DAEB34;
defparam promx9_inst_5.INIT_RAM_27 = 288'h718A1A554AADD72DB6DB6DB6DB6DB75BADD6EB75B6DB6CB5D6683061C11C8A3D32466975;
defparam promx9_inst_5.INIT_RAM_28 = 288'h387B0E7539A3BFDBCD48B4718C30383CA0E371B0EDA4FF7391C6E3B6945C78617D95C6E3;
defparam promx9_inst_5.INIT_RAM_29 = 288'hFBFDF0E845231189AFEB75BADD6DB6DB2B95BAFAF99CCE66A956D10743B9BEDF6737DA71;
defparam promx9_inst_5.INIT_RAM_2A = 288'hEBF5FAFD7EBF5FADB6BAD57AFF7EBD554A84622918987EBF5FEFF7DB31106A4526A3AFF7;
defparam promx9_inst_5.INIT_RAM_2B = 288'hFBFDFEFF7DB75BADD6EB6DBAFD6EB75BADD7EBF5FAFD7EBF5FAFD7FBF5FAFD7EBF5FAFD7;
defparam promx9_inst_5.INIT_RAM_2C = 288'hFBFDFEFF7FBFDFEE17FB85C2E170B85C2FF7FB85C2FF70BFDC2E170BFDFEFF7FBFDFEFF7;
defparam promx9_inst_5.INIT_RAM_2D = 288'hBAF582E17FBFDC2FF70B85FEFF7FB85FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_5.INIT_RAM_2E = 288'hDB6DB6D959A2CB1C48B359ACD66A3516CD467220A4B04A359A8D67082CA19A692614D250;
defparam promx9_inst_5.INIT_RAM_2F = 288'hE73CEEBB6DB75BAFD7EBFDFEFF7FBFDFEFD7EBF5FADD6DB65668928651144827261A08A2;
defparam promx9_inst_5.INIT_RAM_30 = 288'h0701E0903B6BCE2734AA5D72B95CB6DB6DB6DB75BADD6EB75B6DB6CAD51E7CE71B8D44E3;
defparam promx9_inst_5.INIT_RAM_31 = 288'hE6FB7DC6C687B3DBCB7AD4E264C86BC521CD383AD86E361B0C100F2830E4871E738DC786;
defparam promx9_inst_5.INIT_RAM_32 = 288'h82DD7EFD7EBF5ACE843198D498EEB75BADB6DB6DB6B95CA94BD9CBD5EB3598E17349628D;
defparam promx9_inst_5.INIT_RAM_33 = 288'hEBF5FAFD7EBF5FAFD7EBF5AED05633154B06EB75DE905522918946DB75BAFD7FBF5EEAA4;
defparam promx9_inst_5.INIT_RAM_34 = 288'h0BFDFEFF7FBFDFEFF7EB75BADD6EB75BADD7EB75FAFD6EBF5FAFD7EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_5.INIT_RAM_35 = 288'hFBFDFEFF7FBFDFEFF70BFDFEFF7FB85C2FF70BFDFEFF70B85C2E17FBFDFEE170BFDFEE17;
defparam promx9_inst_5.INIT_RAM_36 = 288'h61B0D86C371B8D44AADB05FEE170B85C2FF70BFDFEE17FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_5.INIT_RAM_37 = 288'h5120E0882CAEDB6DB6BACD1658E24E1A8B66B351A8C82A359ACD46A3599868271B8D86C3;
defparam promx9_inst_5.INIT_RAM_38 = 288'h61D95C92538CD32BB6EB75FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFD7EB6DB2B34596B954E3;
defparam promx9_inst_5.INIT_RAM_39 = 288'h71B8DC744F7122480F89C4E27149A552EB95CB65B6DB6DB75BADB6EB6DB6DB6BACD1A4A2;
defparam promx9_inst_5.INIT_RAM_3A = 288'h37CB023126902BDC2C78A2F9BECF6FADE93389344DE71A230D86C371B0ECBCD4881CA0EB;
defparam promx9_inst_5.INIT_RAM_3B = 288'hEBF5EEAC552027AFD7EB7DF5CC44251CE5D6EB75B6DB6DB6572B96CAE57D5ECD5EAF560C;
defparam promx9_inst_5.INIT_RAM_3C = 288'hEBF5FAFD7EB75FAFD7EBF5FAFD7EBF5EAB0572B1588A43975FADD7EB5B948A472B4FEFD7;
defparam promx9_inst_5.INIT_RAM_3D = 288'h0B85FEFF7FBFDFEFF7FBFDFEFF7EB75B6DB6EB75BADD7EB75FAFD6EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_5.INIT_RAM_3E = 288'hFBFDFEFF70B85FEFF7FBFDFEE17FB85FEFF70BFDFEFF70BFDC2E17FB85C2E170BFDC2FF7;
defparam promx9_inst_5.INIT_RAM_3F = 288'h61B0985655130D44A25128D46C371A8925F7FBFDC2FF7FB85FEE17FBFDFEE17FBFDFEFF7;

pROMX9 promx9_inst_6 (
    .DO({promx9_inst_6_dout_w[26:0],promx9_inst_6_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_13),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_6.READ_MODE = 1'b1;
defparam promx9_inst_6.BIT_WIDTH = 9;
defparam promx9_inst_6.RESET_MODE = "SYNC";
defparam promx9_inst_6.INIT_RAM_00 = 288'h9A34B5DA661A0944C38A6DB6DB6DB65668B2D71A70D45A34960966A35164B4651B0D86C3;
defparam promx9_inst_6.INIT_RAM_01 = 288'hBACD1228261A8986E379D532BB6EB75FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5F6D95;
defparam promx9_inst_6.INIT_RAM_02 = 288'h27A430AE371B8DC72307038E33379BCDE734AA5D6EB95CB65B6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_6.INIT_RAM_03 = 288'hE5F3357AB2803B99CB69C49E60A99843DBCCF6FB79BC99A5D164C361B0D86C361B0DC94C;
defparam promx9_inst_6.INIT_RAM_04 = 288'h42292CDB6EBED862A4522920B76DB4B790A4526DBAFB6EB6DB6DB6DB65B2D95CADD669AF;
defparam promx9_inst_6.INIT_RAM_05 = 288'hEB75FAFD7EBF5FAFD7EBF5BADD7EBF5FAFD7EBF5A68C56231188C5932AFADD6DB6DA4AC4;
defparam promx9_inst_6.INIT_RAM_06 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFD7DB6DB6DD6EB75BADD7EBF5BAFD7EBF5FAFD7;
defparam promx9_inst_6.INIT_RAM_07 = 288'hFBFDFEFF70BFDFEFF7FB85FEFF7FBFDFEFF70BFDC2E17FBFDFEFF7FB85FEE170BFDC2E17;
defparam promx9_inst_6.INIT_RAM_08 = 288'h71B8D86A2A2B2CD2C35128944A251A8D47E761B0D86C39A7DFEFF7FBFDFEFF7FB85FEFF7;
defparam promx9_inst_6.INIT_RAM_09 = 288'hFBF5FADB6BACD0A32C40A8A48E3416DBADD6EB6DB2B34596B8936692D168D45A2D168C61;
defparam promx9_inst_6.INIT_RAM_0A = 288'hDB6DB6D96BACD05F245128945E779DD76DB6EB75FAFF7EBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_6.INIT_RAM_0B = 288'h61B0F0D6C58D95C6E371B8DC704D6B4A26F389BCDE734AA556EB75CB6DB6DB6DB6DB6DB6;
defparam promx9_inst_6.INIT_RAM_0C = 288'hAACD1E8D36943757AB8683F95CCE6F2A693389243D9CDE6F379BCE05C4D62C36130D86C3;
defparam promx9_inst_6.INIT_RAM_0D = 288'hDB75E68A452291088472B158AA441A9106836231188A3837DFADD6DB6DB6D96CB5DAEB75;
defparam promx9_inst_6.INIT_RAM_0E = 288'hEB75FAFD7DB75FAFD6EBF5FAFD7EBF5FADD7EBF5FAFD7EBF5B6D8F72B1588C4522914967;
defparam promx9_inst_6.INIT_RAM_0F = 288'hFB85C2E17FBFDC2FF70B85C2FF7FBFDFEFF7FBFDFEFF7DB75BADD6EB75BADD7EBF5BAFD7;
defparam promx9_inst_6.INIT_RAM_10 = 288'hFBFDC2FF7FBFDC2FF7FBFDFEFF7FBFDFEFF7FBFDFEE170BFDFEFF7FB85C2FF70B85C2FF7;
defparam promx9_inst_6.INIT_RAM_11 = 288'h82B0CC4C361A8D5449A230D44A261B0D86C361B0D44A25128946C371A2BEFF7FBFDFEFF7;
defparam promx9_inst_6.INIT_RAM_12 = 288'hFBFDFEFF7FBFDFAFB6CAD51658E4120904A2415D76DD6EB75F6D759A2CB9C48B35168B05;
defparam promx9_inst_6.INIT_RAM_13 = 288'hDB6DB6DB6DB6DB6DB6BACD0A0EB30B8E08C3D75D76DB6EB75FAFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_6.INIT_RAM_14 = 288'h61B0D86C37181C9EB128411C6C371B8DC74C89CD226F389C526934AA5D6EB95CB65B6DB6;
defparam promx9_inst_6.INIT_RAM_15 = 288'hCADD6EB559A451E6D359349628BE50BD9BCCE67B799EBAACCCD9CEF6FB79BCDF644DA2C2;
defparam promx9_inst_6.INIT_RAM_16 = 288'h62B11068431A120AC56231148845231188A45229148836229108A3D3F5BADB6DB6DB6D96;
defparam promx9_inst_6.INIT_RAM_17 = 288'hEB75BAFD6EBF5FADD7EBF5BAFD7EBF5BADD7EBF5FAFD7EBF5FADD6EB75BADF7EBF5B6C4A;
defparam promx9_inst_6.INIT_RAM_18 = 288'hFBFDC2FF7FBFDFEFF7FB85FEFF70B85FEFF7FB85FEFF7FBFDFEFF7DB75B6DD6EBF5FADD7;
defparam promx9_inst_6.INIT_RAM_19 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEFF7FB85FEFF7FB85FEFF7;
defparam promx9_inst_6.INIT_RAM_1A = 288'h1451506E35130A08A361A8986A25130D86C361B0D86C361B0D86C361A8944A25138E49D7;
defparam promx9_inst_6.INIT_RAM_1B = 288'hFBFDFEFF7FBFDFEFF7FBF5FAFB6DB555A56D822898682C75576DD6EBF5FADB6BAC51658D;
defparam promx9_inst_6.INIT_RAM_1C = 288'hCB65B6DB6DB6DB6DD6DB6DB6D95BAD5124EB30B0E08A2045532DB6DB75FAFD7FBFDFEFF7;
defparam promx9_inst_6.INIT_RAM_1D = 288'hF6BD1E58561B0D86E3E69C08E680779DC6E361C13DF139A45227138A4D26954AADD72B95;
defparam promx9_inst_6.INIT_RAM_1E = 288'hDB6DB2D95BADD6AB559A451E6D3692C966B248FBB5DCCE67339BEDF644DE4B1E5F339BCC;
defparam promx9_inst_6.INIT_RAM_1F = 288'hDBEDBAFD6AAB95CAC45231188C55229148A45229148A441A91488341A0D08A4A6EDB6DB6;
defparam promx9_inst_6.INIT_RAM_20 = 288'hEB6DBADD7EBF5FAFD7EBF5FAFD7EBF5BADD6EB75FADD7EBF5FADD7EBF5FADD7EBF5FAFD7;
defparam promx9_inst_6.INIT_RAM_21 = 288'h0B85FEFF7FBFDC2FF70BFDFEFF70BFDC2FF70B85FEFF7FB85C2FF7FBFDFEFF7DB75BADD6;
defparam promx9_inst_6.INIT_RAM_22 = 288'h5130DC744EBFDFEFF7FBFDFEFF7FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEFF7FB85FEE17;
defparam promx9_inst_6.INIT_RAM_23 = 288'hCB555E691A601FCEAA5120986C35128944C361B0D86C361B0D86C361B0D86C361B0D44A2;
defparam promx9_inst_6.INIT_RAM_24 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FADB6CB555A56D5138E8B0475DD76DD6EBF5FADB6;
defparam promx9_inst_6.INIT_RAM_25 = 288'hBADD72B95CB6DB6DB6DB6DB6DB6DB6DB6DB6CADD5E78D61A0904A261FBF6DB6DB75BAFD7;
defparam promx9_inst_6.INIT_RAM_26 = 288'h8984799EDE65BDE50B71B0ECA4F4840DC765D6BADC6E3B294226F379C4DE7138A4D26954;
defparam promx9_inst_6.INIT_RAM_27 = 288'h69EDB6DB6DB65B2B75BAD56AB349A45228F369B4D64B269BCDA44BE67B399ECF6945A52D;
defparam promx9_inst_6.INIT_RAM_28 = 288'hEBF5FAFD7EBF5FAFD7EB6DB50C56231588C46231148A45229148A45228D46A351A0D46A4;
defparam promx9_inst_6.INIT_RAM_29 = 288'hDB6DBADD6EB6DBADD6EB75BADD6EBF5FAFD7EBF5BADD6EB75FADD6EB75BADD6EBF5FAFD7;
defparam promx9_inst_6.INIT_RAM_2A = 288'hFB85C2E170BFDFEFF7FBFDFEFF7FBFDFEE170BFDFEFF70B85C2E170BFDFEFF7FBFDFEFF7;
defparam promx9_inst_6.INIT_RAM_2B = 288'h61B0D86A25161A08E365F5FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_6.INIT_RAM_2C = 288'hEBF5FAFD6DB5D668D2284B206075130D86C35128946C361B0D86C361B0D86C361B0D86C3;
defparam promx9_inst_6.INIT_RAM_2D = 288'hDB75BAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5FADB6BACD165E730A0A48A2145D76DD7;
defparam promx9_inst_6.INIT_RAM_2E = 288'h9A4D2A955BAE572B96CB6DB6DB6DB6DB6DB6DB6DB6DB6CB5D6663065D14C30461A8A69B6;
defparam promx9_inst_6.INIT_RAM_2F = 288'hF6AB5E66CF6F41A4EEE6132263071A249E0F6138DC703D6DB5C62848BCDA6D379C4E2714;
defparam promx9_inst_6.INIT_RAM_30 = 288'h522914745964332D96CB65AEB75AAD56AB349A45228F379B4DA6D369BCDE71328FAFDBED;
defparam promx9_inst_6.INIT_RAM_31 = 288'hEBF5BAFD6EB75BAFD7EBF5FAFD7DBF5FAD1462B1588C46231148A45229148834229148A3;
defparam promx9_inst_6.INIT_RAM_32 = 288'hFBFDFEFF7DB6DB6DB6EB75BADD6EB75FADD6EBF5FADD7EBF5BADD7EBF5BADD7EB75FADD7;
defparam promx9_inst_6.INIT_RAM_33 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF70B85C2E170BFDFEE170B85FEFF7FBFDFEFF70BFDC2FF7;
defparam promx9_inst_6.INIT_RAM_34 = 288'h61B0D86C361B0D86A25128944C351557AFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_6.INIT_RAM_35 = 288'h79DD76DD6EBF5FAFD6DB656A8F348FBDD8074120946A35128D86C361B0D86C361B0D86C3;
defparam promx9_inst_6.INIT_RAM_36 = 288'h411856575DB75BAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5F6D959A14504A261B0D8504;
defparam promx9_inst_6.INIT_RAM_37 = 288'h79C4E29349A552A975BAE572B96DB6DB6DB6DB75BADB6DB75B6DB6DB656A8D3F7C110461;
defparam promx9_inst_6.INIT_RAM_38 = 288'h79C5063CBF68322410F6FB7D6726892A28D10724256E371B8DC6E3E76BA58F279B4DA6F3;
defparam promx9_inst_6.INIT_RAM_39 = 288'h21988C4835130D46A3618A0A396CB5D6EB55AAD5669349A45228F379BCDE6D369BCDE6F3;
defparam promx9_inst_6.INIT_RAM_3A = 288'hEB75BAFD7EB75BAFD6EB75FAFD7EBF5FAFD7EBF5F6FD7DB61D4AE572D1A4AC441A0D0683;
defparam promx9_inst_6.INIT_RAM_3B = 288'h0BFDFEFF7FBFDFEFF7DB75B6DD6DB75BAFD6EB75FAFD6EBF5BADD7EBF5FADD6EBF5BADD7;
defparam promx9_inst_6.INIT_RAM_3C = 288'hFB85FEFF7FBFDFEFF70BFDFEFF70BFDC2FF7FB85C2E170BFDFEFF70B85FEE170BFDC2E17;
defparam promx9_inst_6.INIT_RAM_3D = 288'h61B0D86C361B0D86C361B0D86C361A8944A261823ADD7EBFDFEFF7FBFDFEFF7FB85C2FF7;
defparam promx9_inst_6.INIT_RAM_3E = 288'h82208D2309A6576DD7EBF5FAFD6DB656A913488BE18E441209C8E45128D86A351B0D86C3;
defparam promx9_inst_6.INIT_RAM_3F = 288'h38BAD84615138D8628CAEDBADD7FBFDFEFF7FBFDFEFF7FBFDFEFF7EB6DB2D5579C90C504;

pROMX9 promx9_inst_7 (
    .DO({promx9_inst_7_dout_w[26:0],promx9_inst_7_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_15),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_7.READ_MODE = 1'b1;
defparam promx9_inst_7.BIT_WIDTH = 9;
defparam promx9_inst_7.RESET_MODE = "SYNC";
defparam promx9_inst_7.INIT_RAM_00 = 288'h79BCDE6F38A4D26934AA556AB75BAE572DB6CB6DB6DB6DB75BADD6EB75BADB6DB656EB34;
defparam promx9_inst_7.INIT_RAM_01 = 288'h79BCDE6F379BCE2913F8F322891077B79A0EF5ACA22D278F9D86E371B8DC6E307F3A2713;
defparam promx9_inst_7.INIT_RAM_02 = 288'h3198D88E562188C48340A0904623120ACB75BADD6AB55AACD269149A452291479BCDE6F3;
defparam promx9_inst_7.INIT_RAM_03 = 288'hEBF5FADD6EB75BAFD6EB75BAFD6DB75FAFD7EBF5FAFB6EBF5FAFD7EBF5FADB6EB24A4AC3;
defparam promx9_inst_7.INIT_RAM_04 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7DB6DBADD6DB75BADD6EB75FADD7EB75BADD7EBF5FADD6;
defparam promx9_inst_7.INIT_RAM_05 = 288'hFBFDFEFF7FBFDFEE17FB85C2E17FB85FEFF70B85FEFF70BFDFEE170B85C2E17FB85C2E17;
defparam promx9_inst_7.INIT_RAM_06 = 288'h61B0D86C361B0D86C361B0D86C35128986C361A89442861A8B6DD6EBFDFEFF7FBFDFEFF7;
defparam promx9_inst_7.INIT_RAM_07 = 288'h6138D444161A082113CAEDBADD7EBF5FAFD6DB656A8F33883C90C35120946A35128D86C3;
defparam promx9_inst_7.INIT_RAM_08 = 288'hDB6DB2B5479FBD55244169ECCC38A6DB6DD6EBF5FAFF7FBFDFEFF7EBF5FADD6DB656A8D2;
defparam promx9_inst_7.INIT_RAM_09 = 288'h2844E26F379BCE27139A4D26954AAD56EB75CAE5B2DB6DB6DB6DB6DB6DBADD6EB75BADB6;
defparam promx9_inst_7.INIT_RAM_0A = 288'h8A3CDE6F379C5229148A3CDE71389C5120B2F67B7D9CDF6737D5122830D86E371B0DC765;
defparam promx9_inst_7.INIT_RAM_0B = 288'hDB491C8C361A90C6634229106614120944A3412094786AAD5669349A4D269148A4522914;
defparam promx9_inst_7.INIT_RAM_0C = 288'hEBF5BADD7EB75FADD6EBF5BADD7EB75B6DB6EB75BAFD7EBF5FAFD7EBF5FAFD7DBEDB6DB6;
defparam promx9_inst_7.INIT_RAM_0D = 288'hFBFDC2E170B85FEFF7FBFDFEFF7FBFDFEFF7DB6DB6DD6EB6DBADD6EB6DBADD6EB75BAFD6;
defparam promx9_inst_7.INIT_RAM_0E = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2FF7FBFDC2E17FBFDFEFF7FBFDC2FF70B85C2E17;
defparam promx9_inst_7.INIT_RAM_0F = 288'h51A8986C361B0D86C361B0D86C351A8D46A35128D46C361A8944A251A8A27D6EBF5FEFF7;
defparam promx9_inst_7.INIT_RAM_10 = 288'hBABCDA4A271D9A088271CB1A555DB75BADD7EBF5FADD6DB65AA8F338FBECB255128986C3;
defparam promx9_inst_7.INIT_RAM_11 = 288'hEB75BADB6DB6DB2D759A2CB9D24412898661595D76DB6EB75FAFD7EBF5FAFD7EBEDB6D96;
defparam promx9_inst_7.INIT_RAM_12 = 288'h61B0FCE7089C4DE6F389C4E29349A552A955AAD56EB75CAE5B2DB6DB6DB6DB6DB6DBADD6;
defparam promx9_inst_7.INIT_RAM_13 = 288'h8A45229148A45229148A45229148A45229148A4D2A934C7FB3D9ECE6733DAF258B8D86C3;
defparam promx9_inst_7.INIT_RAM_14 = 288'hEBF5FAFB60838DC6825120906A44198544824120904A3512090504F7CD269148A4522914;
defparam promx9_inst_7.INIT_RAM_15 = 288'hEB75FAFD7EBF5BAFD6EB75BADD6EB75BAFD6DB75FADB6EB75BAFD7EBF5FAFD7EBF5FAFB6;
defparam promx9_inst_7.INIT_RAM_16 = 288'h0BFDFEFF7FBFDC2E170BFDFEE17FB85FEFF7FBFDFEFF7DB75B6DB6DB6DBADD6DB6DBADD7;
defparam promx9_inst_7.INIT_RAM_17 = 288'hEB75FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2FF7FBFDC2FF7;
defparam promx9_inst_7.INIT_RAM_18 = 288'h5130944C361A8944C361B0D86C361B0D86C351B0D46A351A8D46C35128944A261A8965D6;
defparam promx9_inst_7.INIT_RAM_19 = 288'hDB656A96D61A89046141209C882D734AAB96DB75FAFD7EBF5FAFD6DB65AEB1338F3810A3;
defparam promx9_inst_7.INIT_RAM_1A = 288'hDB75B6DD6EB75BADD6EB6DB6D96BAC4CA0EB7210546E361EBB2BB6DB75BADD6EB75BADD6;
defparam promx9_inst_7.INIT_RAM_1B = 288'h6830986C371AA962F379BCDE71389C5269349A552AB55BADD6EB95CAE5B6DB6DB6DB6DB6;
defparam promx9_inst_7.INIT_RAM_1C = 288'h79BCE29148A45229148A45269349A4D269349A4D269349A4D269549A34817CCE6733DBF0;
defparam promx9_inst_7.INIT_RAM_1D = 288'hDB6DB6DB6DB6DB6DB61430D86E351A0DC8E351209C8C37239186C361A0904A21445228F3;
defparam promx9_inst_7.INIT_RAM_1E = 288'hEB75BADD6EB75BAFD7EB75FADD7EB75BADD6EB75BADD6EB75BADD6EB75BAFD7DB75FAFD7;
defparam promx9_inst_7.INIT_RAM_1F = 288'h0B85C2FF70B85C2FF70B85C2FF7FBFDC2FF7FBFDFEFF7FBFDFEFF7DB6DB6DD6EB75B6DD6;
defparam promx9_inst_7.INIT_RAM_20 = 288'h51209A7B6EB75FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70BFDC2FF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_7.INIT_RAM_21 = 288'h59739D76551289C6A261B0D44A261B0D86C361B0D86C361B0D86A351A8D44C361A8944C2;
defparam promx9_inst_7.INIT_RAM_22 = 288'hDB6DAEB75C730FCE8261C91864130A89C90B695576DB6EBF5FEFF7EBF5FAFD6DB656EB34;
defparam promx9_inst_7.INIT_RAM_23 = 288'hDB6DB6DB6DB75BADD6EB75BADD6EB75B6DB6BAD51A5CF4530987A792B0E6995CAE5B6DB6;
defparam promx9_inst_7.INIT_RAM_24 = 288'hF5F33DA8C7881DC6E3C6B49E6D279C4E27148A4D26954AAD52AB75BADD6EB95CAE5B6DB6;
defparam promx9_inst_7.INIT_RAM_25 = 288'hD33ADA6D379B4DE6F379C5229148A4D269349A4D269349A4D269349A4D269148A3CE2693;
defparam promx9_inst_7.INIT_RAM_26 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6D9671A8D86E371B92092592A8E094592C11C8E361A890482;
defparam promx9_inst_7.INIT_RAM_27 = 288'hEB75BADD6EB75BADD6EBF5BADD6DB75BADD6EB75BADD6EBF5BADD6EB75BADD6EB75B6DD7;
defparam promx9_inst_7.INIT_RAM_28 = 288'h0BFDC2E17FBFDC2E170B85C2FF7FBFDFEFF70C05FEFF7FBFDFEFF7FBFDFEFF7DB75BADB6;
defparam promx9_inst_7.INIT_RAM_29 = 288'h5128944A372412AB96DB75BAFD7EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_7.INIT_RAM_2A = 288'hEB6DB2B54798C2586971A09C6C35130D86A25130D86C361B0D86C361B0D86A351A8944A2;
defparam promx9_inst_7.INIT_RAM_2B = 288'h71E1AAB551438D65864130D44822098504C3142271CB2AA65B6DD6EBFDFEFF7FBFDFAFD7;
defparam promx9_inst_7.INIT_RAM_2C = 288'hCB6DB6DB6DB6DB6DB6EB75BADD6EB75BADD7EBF5B6DB6CADD668B2E730D44C3A290596A2;
defparam promx9_inst_7.INIT_RAM_2D = 288'h8A451E6F3798C797EB796B289EF89BCDE6F379C4E69349A4D2A955AAD56EB75CAE572B96;
defparam promx9_inst_7.INIT_RAM_2E = 288'h61A0944C3B2F1D64B25934DA6F379C5229149A4D269349ACD66B55AAD56AB559A4D26934;
defparam promx9_inst_7.INIT_RAM_2F = 288'hEB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB2D96D328D86E4724128B46A3391472592C11C6C3;
defparam promx9_inst_7.INIT_RAM_30 = 288'hDB6DB6DB6EB6DBADD6EB75BADD7EBF5BAFD7EB75B6DD6EB75BADD6EB6DBADD6EB75BADD6;
defparam promx9_inst_7.INIT_RAM_31 = 288'h0BFDFEFF7FB85FEE170B85FEE17FB85C2FF7FB85FEE17FB85FEE170BFDFEFF7FBFDFAFF7;
defparam promx9_inst_7.INIT_RAM_32 = 288'h5128944A251A8946C34138EEBB6DB75BAFD7FBFDFEFF7FBFDFEFF7FBFDFEE17FBFDFEE17;
defparam promx9_inst_7.INIT_RAM_33 = 288'hFBFDFAFD7EB6DB2B5489ACB9CEA1428944E361A8986C35128944C361B0D86C361A8986A3;
defparam promx9_inst_7.INIT_RAM_34 = 288'h4130CC4E3A2C10C2615130D46414120986614130E078D2834A2775DB75BADF7FBFDFEFF7;
defparam promx9_inst_7.INIT_RAM_35 = 288'hCAE572D96DB6DB6DB6DB6DB6DB6EB75BADD6EB75BADD6EB75BADB6DB656AB130879DC6A2;
defparam promx9_inst_7.INIT_RAM_36 = 288'hAAD56AB559A4D228F379BCDE610792C4E13389C4E27138A4D26954AA556AB55BADD6EB75;
defparam promx9_inst_7.INIT_RAM_37 = 288'h51A0944A24128944C3A29A52492592C964D379C5229349A4D6AB35AAD56AB55AAD56AB55;
defparam promx9_inst_7.INIT_RAM_38 = 288'hEB75BADD6DB6DBADB6DB6DB6DB6DB6DB6DB6DB65B2D96C739186E4724168B45A2B910504;
defparam promx9_inst_7.INIT_RAM_39 = 288'hFBFDFEFF7DB6DB6DB6DB6DBAFB6EB75BADD6EB75FADD6EB75BAFD7EB75BADD6EB6DBADD6;
defparam promx9_inst_7.INIT_RAM_3A = 288'hFBFDFEFF7FBFDFEFF7FB85FEFF70B85FEFF70B85FEFF7FB85FEE17FB85FEFF7FBFDFEFF7;
defparam promx9_inst_7.INIT_RAM_3B = 288'h61A8944A25128944A261A8D46A3E3F1B2B96DB75BAFF7FBFDFEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_7.INIT_RAM_3C = 288'hFBFDFEFF7FBFDFEFF7EB75B6D759A3CCE3AE650A102A261B0D44C371B0F4CE35130D86C3;
defparam promx9_inst_7.INIT_RAM_3D = 288'h6973955C7C369904C361B0CC2614130D44CA40989054575D341ED29A5D72DB6EBFDFEFF7;
defparam promx9_inst_7.INIT_RAM_3E = 288'hBADD72B95CAE5B2DB6DB6DB6DB6DB75BADB6EB75BADD6EB75BADD6EBF5FADB6DB6DB2B54;
defparam promx9_inst_7.INIT_RAM_3F = 288'hBADD6EB55AAD56AB55AACD269149A4D26B75CAEDB2B559A4D269349A4D2A955AAD56EB75;

pROMX9 promx9_inst_8 (
    .DO({promx9_inst_8_dout_w[26:0],promx9_inst_8_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_17),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_8.READ_MODE = 1'b1;
defparam promx9_inst_8.BIT_WIDTH = 9;
defparam promx9_inst_8.RESET_MODE = "SYNC";
defparam promx9_inst_8.INIT_RAM_00 = 288'h51A8904A24120904825120986E4548C0A271492C964D379C5229349A556AB55AAD56AB55;
defparam promx9_inst_8.INIT_RAM_01 = 288'hEB6DBADB6EB75BADB6EB6DB6DB6DB6DB6DB6DB6DB6D96CB65B2D969A69944A3624968CE4;
defparam promx9_inst_8.INIT_RAM_02 = 288'hFBFDFEFF7FBFDFEFD7DB6DB6DD6DB75FAFD6EB75BADD7EBF5BADD6EBF5BADD7EB75B6DD6;
defparam promx9_inst_8.INIT_RAM_03 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FB85FEFF7FBFDC2FF70B85C2FF7FBFDC2FF7FBFDFEFF7;
defparam promx9_inst_8.INIT_RAM_04 = 288'h61B0D86A25128944A25128946C361B8DC607925B6EB96DB75BADF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_8.INIT_RAM_05 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5B6D95AA4D1A450C6AA850815120904825130D86E3;
defparam promx9_inst_8.INIT_RAM_06 = 288'hEB6DB6D96BAC4D6450F7BAE06A25130F4CA24120B8F4C34D9513CF5944EA976DB6DBADD7;
defparam promx9_inst_8.INIT_RAM_07 = 288'hBADD6EB75CAE572B95CB65B6DB6DB6DB6DB6EB75B6DD6EB75BADD6EB75FADD7EBF5FAFD6;
defparam promx9_inst_8.INIT_RAM_08 = 288'hAAD56EB75BADD6EB75AAD56AB75BAD56AB55AAD56EB95EB75B2B95AADD6AB55AAD56EB75;
defparam promx9_inst_8.INIT_RAM_09 = 288'h6259ACCE451A0904A24128944A251289C606B503C605138A4964D379C526934AAD56AB55;
defparam promx9_inst_8.INIT_RAM_0A = 288'hEB75BADD6EB75BADD6EB75BADD6DB6DB6DB6DB6DB6DB6DB6DB6DB6CB65B2D75BABAECAC3;
defparam promx9_inst_8.INIT_RAM_0B = 288'hFB85FEFF7FBFDFEFF7FBFDFEFF7EB6DB6DD6DB6DBADD6EB75BADD6EB75FADD6EB75BAFD6;
defparam promx9_inst_8.INIT_RAM_0C = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF70B85FEFF7FBFDFEFF7FBFDFEFF70B85FEFF70B85C2FF7;
defparam promx9_inst_8.INIT_RAM_0D = 288'h61A0904A261B0DC6E361B0D86C361B0D86A34120A8B44820C2EB96DB75BAFD7FBFDFEFF7;
defparam promx9_inst_8.INIT_RAM_0E = 288'hEB75FEFF7FBFDFEFF7FBFDC2E17FBFDFEFF7EBF5F6DB6BAD5266D228635540771A894482;
defparam promx9_inst_8.INIT_RAM_0F = 288'hEBF5FAFD7EB75BADB6DB65AAB34698C2982803B2E5889C3719956CE7141A734BAE5B6DB6;
defparam promx9_inst_8.INIT_RAM_10 = 288'hBADD6EB75BAE572B95CB65B2D96DB6DB6DB6DB6DB6DB6EB75BADD6EB75BADD6EB75FAFD7;
defparam promx9_inst_8.INIT_RAM_11 = 288'h9AD56AB55AADD6EB75BADD6ED76BADD6EB95BADD6EB75BAE5B2DB6DB6DB2D96CADD6EB75;
defparam promx9_inst_8.INIT_RAM_12 = 288'hAAB4C1125824964AE48228904825128944A251B0EC92AB5FBC203028A4964D379C526934;
defparam promx9_inst_8.INIT_RAM_13 = 288'hEB75FADD6EB75BADB6DB75BADB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2D96CB65B2D75;
defparam promx9_inst_8.INIT_RAM_14 = 288'h0B85C2E170BFDFEFF7FBFDFEFF7FBFDFEFF7DB6DB6DD6EB75FADD6EB75BADD6EB75BADD6;
defparam promx9_inst_8.INIT_RAM_15 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2E170BFDC2E170BFDFEE170B85C2E17;
defparam promx9_inst_8.INIT_RAM_16 = 288'h1420986A271A0904A25120986C39241186A241184C26141208C461511C2EB96DB75BAFD7;
defparam promx9_inst_8.INIT_RAM_17 = 288'hDB75BAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FADB6CADD6A913691431ACA;
defparam promx9_inst_8.INIT_RAM_18 = 288'hEBF5BAFD7EBF5FAFD6EBF5FADD6EB6DB6D95BACD1E6B248AC9A49238940A18D58CD2EBB6;
defparam promx9_inst_8.INIT_RAM_19 = 288'hCAE572B95CAE572B95CAE5B2D96CB65B2DB6DB6DB6DB6DB6DB6DD6EB6DBADD6EB75BAFD7;
defparam promx9_inst_8.INIT_RAM_1A = 288'h7A4526935AAD56AB75BADD72B75BAE572B96BAE572B95CAE5B2D96CB6DB6DB6DB6DB6D96;
defparam promx9_inst_8.INIT_RAM_1B = 288'hCB65AEB75AAD57CFA7A2C1208E461A8D44825120902A254B25952BC673FDE3038A4964D3;
defparam promx9_inst_8.INIT_RAM_1C = 288'hEB75BADD7EB75BADD6EB75BADD6EB75BADD6EB75B6DB6EB6DB6DB6DB6DB6DB6DB65B2D96;
defparam promx9_inst_8.INIT_RAM_1D = 288'hFB85C2E170B85C2E17FB85FEFF7FBFDFEFF7FBFDFEFF7DB6DBADB6EB75B6DD6EB75BADD6;
defparam promx9_inst_8.INIT_RAM_1E = 288'hDB75BAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70B85C2E17FB85FEFF70B85FEE17;
defparam promx9_inst_8.INIT_RAM_1F = 288'h89B48E3CE75121C6A25130D868261B0DC70471B0D046230984C26120C128D875171E6996;
defparam promx9_inst_8.INIT_RAM_20 = 288'hBA9C76DD6EBF5FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FAFB6DB656EB54;
defparam promx9_inst_8.INIT_RAM_21 = 288'hEBF5FADD7EB75FAFD7EBF5FAFD7EBF5FAFD7EB75F6DB6DB65AEB75BADD6EB55AAD526954;
defparam promx9_inst_8.INIT_RAM_22 = 288'hDB6DB6DB6CB65B2D96DB6DB2D96CB65B2D96CB6DB6DB6DB6DB6DB6DB6DB6DD6EB75BADD6;
defparam promx9_inst_8.INIT_RAM_23 = 288'h38AC9A4F38A4D2A955AADD6EB75CAE572B95CB6572D95CB65B2D96DB6DB2DB6DB6DB6DB6;
defparam promx9_inst_8.INIT_RAM_24 = 288'hDB6DB2D96CB65AEB75AAD566914F7D12490571B0D86C2E2CAA554AA5529112BC6EB81E50;
defparam promx9_inst_8.INIT_RAM_25 = 288'hEB75BAFD6EBF5BAFD6EB75BADD6EB75BADD6DB75BADD6EB75BADB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_8.INIT_RAM_26 = 288'hFBFDFEFF7FB85FEE170BFDC2E17FBFDC2FF70B85FEFF7FBFDFEFF7DB6DBADB6EB75BADD6;
defparam promx9_inst_8.INIT_RAM_27 = 288'hB359F4F54EB75BADD7FBFDFEFF7FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEE17FB85C2FF7;
defparam promx9_inst_8.INIT_RAM_28 = 288'hEB6DB2B75AA44DE671F7D3155A661289C6A28241208E371A08C26131188C505A359ACD66;
defparam promx9_inst_8.INIT_RAM_29 = 288'hDB6572B95CAEDBADD7EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2FF7FBFDFEFF7FBFDFAFD7;
defparam promx9_inst_8.INIT_RAM_2A = 288'hEB75BADD6EBF5FADD7EBF5FAFD6EBF5FAFD7EBF5FEFD7EBF5FAFD6EB75BADB6DB6DB6DB6;
defparam promx9_inst_8.INIT_RAM_2B = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2DB6DB6DB6DB6DB6DB6DB6EB75BADB6;
defparam promx9_inst_8.INIT_RAM_2C = 288'hB6EB8607148B49E7139A4D2A955AADD6EB95CAE5B2B96CB65B2D96CB65B6DB6DB6DB6DB6;
defparam promx9_inst_8.INIT_RAM_2D = 288'hDB6DB6DB6CB6DB2D96CB5D6EB75BAD56691479B409DCC44EB3158AC562B156AC5E30914C;
defparam promx9_inst_8.INIT_RAM_2E = 288'hEB75B6DD6EB75BADD6EB75BADD6DB75BADD6EB75BADD6EB75B6DD6EB6DBADD6DB6DB6DB6;
defparam promx9_inst_8.INIT_RAM_2F = 288'hFB85C2FF7FB85C2E17FB85C2E170BFDC2E17FBFDFEFF7FB85FEFF7FBFDFEFF7EB6DB6DD6;
defparam promx9_inst_8.INIT_RAM_30 = 288'hB359A8F67B3E1ECDE8CB6DBADD7EBFDFEFF7FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_8.INIT_RAM_31 = 288'hFBFDFEFF7EB75B6D95BAD5268F3590C35D2C75A24938571B8D86E371B0CC4816251A8D46;
defparam promx9_inst_8.INIT_RAM_32 = 288'hEB75BADD6DB6DB6DB6EB75BAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2E17FBFDFEFF7;
defparam promx9_inst_8.INIT_RAM_33 = 288'hDB75BADD6EB75BADD6EBF5FADD7EBF5FAFF7EBF5FAFD7EBF5FAFD7FBF5FAFF7EBF5FAFD6;
defparam promx9_inst_8.INIT_RAM_34 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6CB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_8.INIT_RAM_35 = 288'hA31B1592CC6840A07159349E7149A552AB75BADD72B95CB65B2D96CB6DB6DB6CB6DB6DB6;
defparam promx9_inst_8.INIT_RAM_36 = 288'hDB6DB6DB6DB6DB6DB6DB65B2D96CB65AEB75BAD5669338A3CD627044AA3D9CBE5E2E55C6;
defparam promx9_inst_8.INIT_RAM_37 = 288'hDB6DB6DB6EB6DBADD6EB75FADD6EB75BADD6EB75BADD6EB75BADB6EB75BADD6EB6DB6DD6;
defparam promx9_inst_8.INIT_RAM_38 = 288'hFBFDFEE170BFDFEFF7FBFDC2FF70BFDC2E170B85FEFF7FB85C2FF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_8.INIT_RAM_39 = 288'hA359ACD66B3D9B0D6751C970F87256DBAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_8.INIT_RAM_3A = 288'hFBFDFEFF7FBFDFEFF7FBF5FADB6DB656EB549A3CD64711873B5D6D862AF0CC334F1CC241;
defparam promx9_inst_8.INIT_RAM_3B = 288'hFBFDFAFD7EBF5FAFD7EBF5BADD7EB7DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_8.INIT_RAM_3C = 288'hDB6DB6DD6EB75BADD6EB75BAFD6EBF5FADD6EBF5FAFD7EBF5FAFD7EBFDFAFF7FBFDFEFF7;
defparam promx9_inst_8.INIT_RAM_3D = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6;
defparam promx9_inst_8.INIT_RAM_3E = 288'h7712F0D25A3A2E1B2C0794122B269BCE29349A556EB75BADD72B96CB65B2D96CB6DB6DB6;
defparam promx9_inst_8.INIT_RAM_3F = 288'hEB6DB6DD6EB75B6DB6DB6DB6DB6CB65B2D96CB65AEB75BAD56A9349A3CDE6D248943CB25;

pROMX9 promx9_inst_9 (
    .DO({promx9_inst_9_dout_w[26:0],promx9_inst_9_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_19),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_9.READ_MODE = 1'b1;
defparam promx9_inst_9.BIT_WIDTH = 9;
defparam promx9_inst_9.RESET_MODE = "SYNC";
defparam promx9_inst_9.INIT_RAM_00 = 288'hFBFDFEFF7DB6DB6DD6EB75B6DD6EB75BADD6EB75BAFD7EB75BADD6EB75BADD6EB75BADB6;
defparam promx9_inst_9.INIT_RAM_01 = 288'hFBFDFEE17FBFDFEFF70B85FEFF7FBFDC2E170BFDFEFF7FBFDFEFF7FBFDC2E170B85FEFF7;
defparam promx9_inst_9.INIT_RAM_02 = 288'h921A48387B351ACD66B361CC4E4C3D9B0F87D3AAF6DD6FBFDFEFF7FBFDFEFF7FBFDC2FF7;
defparam promx9_inst_9.INIT_RAM_03 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAFD6DB6DB2D95BAD52691379AC96471288435C28;
defparam promx9_inst_9.INIT_RAM_04 = 288'hEBF5FAFD7EBF5FAFD7FBFDFEFF7EBF5FAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_9.INIT_RAM_05 = 288'hDB6DB6DB6EB6DBADD6EB75BADD6EB75BADD7EB75FADD7EBF5FAFD7EBF5FAFD7EBFDFAFD7;
defparam promx9_inst_9.INIT_RAM_06 = 288'hDB6DB6DB6DB6DB6DB6DB6DBADB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_07 = 288'h591C45123723B65F4FF822AD80F2824564D379C526954AADD6EB95CAE572D96CB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_08 = 288'hEB6DBADD6EB75BADB6EB6DB6DB6DB6DB6DB6DB65B2D96CB65B2D96BAD56A9549A451E6F3;
defparam promx9_inst_9.INIT_RAM_09 = 288'hFBFDFEFF7FBFDFEFF7DB6DBADB6EB6DBADD6EB75BADD6EBF5BADD6EB75BADD6EB75BADD6;
defparam promx9_inst_9.INIT_RAM_0A = 288'hFBFDFEE17FBFDC2FF7FBFDFEFF70B85FEFF70BFDFEE17FBFDC2E170B85C2E17FB85FEFF7;
defparam promx9_inst_9.INIT_RAM_0B = 288'h79AC8E3EF44C968B46C359F0D8630D194621B3E1A0966A361E19B6EBF5FEFF7FBFDFEFF7;
defparam promx9_inst_9.INIT_RAM_0C = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFD7EB6DB6DB6CB656EB55AA4D228F3;
defparam promx9_inst_9.INIT_RAM_0D = 288'hEBFDFAFD7EBF5FAFD7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_9.INIT_RAM_0E = 288'hDB6DB6DD6EB75B6DD6EB75BADD6EB75BADD6EB75BAFD7EB75BAFD7EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_9.INIT_RAM_0F = 288'hCB65B6DB6DB6DB6DB6DB6DB6DB6DB75B6DD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_10 = 288'hAA4D2691379B48A089E301DD74DC703CE29159349E6F38A4D26955BADD6EB95CB6572B96;
defparam promx9_inst_9.INIT_RAM_11 = 288'hEB75BADD6DB6DBADD6DB6DBADB6DB6DB6DB6DB6DB6DB6DB6DB6D96CB65B2B95BADD6EB55;
defparam promx9_inst_9.INIT_RAM_12 = 288'hFB85C2FF7FBFDFEFF7FBFDFEFF7DB6DB6DB6DB75BADD6EB75BADD6EB75BADD6EBF5BAFD6;
defparam promx9_inst_9.INIT_RAM_13 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70BFDFEFF7FBFDFEFF70BFDC2E170BFDFEE17;
defparam promx9_inst_9.INIT_RAM_14 = 288'hCADD6EB559A44E26D22842F0D46B361C8367D3D9F0F6741C970F25C3E1F0F2DEB75FAFF7;
defparam promx9_inst_9.INIT_RAM_15 = 288'hEBF5BADD6CB75B6DF7FBFDFEE17FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5FADB6DB6DB6B95;
defparam promx9_inst_9.INIT_RAM_16 = 288'hEBF5FAFD7EBF5FAFF7EBF5FAFD7EBF5FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FEFD7;
defparam promx9_inst_9.INIT_RAM_17 = 288'hDB6DB6DB6DB6DB6DD6EB75BADD6EB75BADD7EB75BADD6EB75BADD7EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_9.INIT_RAM_18 = 288'hCB6572B95CB65B6DB6DB6DB6DB6DB6DBADB6DB75BADD6EB6DB6DB6DB6DB6DB6DB6DB6D96;
defparam promx9_inst_9.INIT_RAM_19 = 288'hCADD6EB75BAD52A93489BCDA4B248940E2B159349A4D379BCE29349A552A975BADD72B95;
defparam promx9_inst_9.INIT_RAM_1A = 288'hEB75BADD6EB75B6DD6EB6DB6DB6EB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB65B2D95;
defparam promx9_inst_9.INIT_RAM_1B = 288'h0B85C2E17FBFDFEE17FBFDFEFF7FBFDFEFF7DB6DB6DD6DB6DBADD6EB75BADD6EB75BAFD6;
defparam promx9_inst_9.INIT_RAM_1C = 288'hB6E5BAFF7FBFDFEFF7FBFDC2E170BFDFEFF7FBFDFEFF7FBFDC2FF7FBFDFEE17FBFDFEFF7;
defparam promx9_inst_9.INIT_RAM_1D = 288'hEBEDB6DB6DB6DB2B95CADD6A934799C61986A359B0F87C361D0586310830F66B3E1E0B67;
defparam promx9_inst_9.INIT_RAM_1E = 288'hEBF5F6D5407EBB0AC35130DC7B6EBFDFEFF7FBFDFEFF70BFDFEFF7FBFDFEFF7FBFDFAFD7;
defparam promx9_inst_9.INIT_RAM_1F = 288'hEBF5FAFD7EBF5FAFD7EBFDFAFD7FBF5FAFD7FBF5FEFF7EBF5FAFD7EBFDFAFD7FBFDFAFD7;
defparam promx9_inst_9.INIT_RAM_20 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DD6EB75BADD6EB75BADD6EB75FAFD6EB75BAFD6EBF5FAFD7;
defparam promx9_inst_9.INIT_RAM_21 = 288'hBAE572B95BADD72B95CAE572DB6DB6DB6DB6EB75BADD6EB6DB6DB6DB75BADD6DB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_22 = 288'hDB6DB2D95CB6572B75BADD6AB54AA4D2671379BCDE6F379BCDE6F38A4D26954AA556EB75;
defparam promx9_inst_9.INIT_RAM_23 = 288'hEB75BAFD6EB75BADD6EB75FADD6EB6DBADD6DB6DB6DD6EB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_24 = 288'hFBFDFEFF70B85C2FF7FB85C2E17FBFDFEE17FBFDFAFF7DB6DB6DB6DB75B6DD6EB75BADD6;
defparam promx9_inst_9.INIT_RAM_25 = 288'hB3392CF87C3DBBAFF7FBFDFEFF7FBFDFEE17FBFDFEFF7FBFDFEFF70BFDFEFF7FB85FEE17;
defparam promx9_inst_9.INIT_RAM_26 = 288'hFBFDFAFD7EBFDFAFD7EBF5BADB6DB6DB2B95AA44CE34CD359B0F8710D9F0D87B3D99C946;
defparam promx9_inst_9.INIT_RAM_27 = 288'hFBFDFAFD6DB5D5A2A35128986E371B8E4996EBFDFEFF7FBFDC2FF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_9.INIT_RAM_28 = 288'hEB75BAFD7EBF5FAFD7EBF5FAFD7EBFDFAFD7EBFDFEFF7EBF5FAFD7EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_9.INIT_RAM_29 = 288'hEB6DB6DB6DB6DB6DB6DB6DB6DB6DB75B6DD6EB75BADD6EB75BAFD6EB75FAFD6EBF5BADD7;
defparam promx9_inst_9.INIT_RAM_2A = 288'hAADD72B55BAE56EB75AADD6EB75BAE572DB6DB6DB6DD6EB75BADB6DB75B6DD6EB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_2B = 288'hDB6DB6DB6DB6DB6D96DB65B2D95CADD6EB75AAD52A9349A44E271389C5269349A556AB55;
defparam promx9_inst_9.INIT_RAM_2C = 288'hDB6DBAFD6EB75FADD6EB75BADD6DB75BADD6EB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_2D = 288'h0B85FEFF7FBFDFEE170B85C2E170B85C2FF7FBFDFEFF7FBFDFEFF7DB65B6DB6DB6DB6DD6;
defparam promx9_inst_9.INIT_RAM_2E = 288'h6259CC200B359F4F872159F5FD6FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_9.INIT_RAM_2F = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFD7EBF5BADD6EB75B6DB6CADD628919669ACD67C3E1F0F87;
defparam promx9_inst_9.INIT_RAM_30 = 288'hEBF5BAFD6DB6DB2B6BA4C2718E3718235CD2AA5D76DD7FBFDFEFF7FBFDC2FF7FBFDFEFF7;
defparam promx9_inst_9.INIT_RAM_31 = 288'hEBF5BAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBFDFAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7;
defparam promx9_inst_9.INIT_RAM_32 = 288'hEB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6DB75B6DD6EB75FADD6EB75BADD7EB75FAFD6;
defparam promx9_inst_9.INIT_RAM_33 = 288'hAA556EB75BADD6686151536A954AA556AB55BAE572B96DB6DB6DD6EB75BADD6EB75BADD6;
defparam promx9_inst_9.INIT_RAM_34 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2D96CB6572B95BADD6AB55AAD56A954AA4D2A954;
defparam promx9_inst_9.INIT_RAM_35 = 288'hDB6DBADD6EB75B6DD6EB75FADD6EB75BADD6DB75BADB6EB75B6DB6EB6DB6DB6DB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_36 = 288'hFBFDFEFF7FB85FEE17FBFDFEFF70BFDC2E170B85C2FF7FBFDFEFF7FBFDFEFF7DB6DB6DB6;
defparam promx9_inst_9.INIT_RAM_37 = 288'hD3E1C43876261F0F87B359E4A83B3E1F0FAFEB7DFEFF7FBFDFEE17FBFDC2FF7FB85FEE17;
defparam promx9_inst_9.INIT_RAM_38 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5FAFD6DB65AEB3448D330D66;
defparam promx9_inst_9.INIT_RAM_39 = 288'hEB75FADB6CB6D5A2C9A54275A30694D2AB75BAE5B6DB6EB75BAFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_9.INIT_RAM_3A = 288'hEB75FAFD7EB75FAFD7EB75BAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFD7EBF5FAFF6;
defparam promx9_inst_9.INIT_RAM_3B = 288'hEB75BADD6EB75BADD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6EB75BADD6EB75BADD6;
defparam promx9_inst_9.INIT_RAM_3C = 288'hBADD6EB55BADD6EB75AA9A5854CA2B0D04A2F3CD26954AADD72B96DB6DBADD6EB75BADD6;
defparam promx9_inst_9.INIT_RAM_3D = 288'hDB6DB6DB6DB6DB6DB6EB6DB6DB6DB6DB6DB6DB6DB6DB6DB65B2D96CAE56EB75BADD6EB75;
defparam promx9_inst_9.INIT_RAM_3E = 288'hDB6DB6DB6DB75BADD6EB75B6DD7EB75FADD6DB75BADD6EB6DBADB6DB75BADB6EB75BADB6;
defparam promx9_inst_9.INIT_RAM_3F = 288'hFBFDFEFF70BFDC2FF7FBFDFEE170BFDFEE170B85C2E170B85FEFF7FBFDFEFF7FBFDFEFF7;

pROMX9 promx9_inst_10 (
    .DO({promx9_inst_10_dout_w[26:0],promx9_inst_10_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_21),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_10.READ_MODE = 1'b1;
defparam promx9_inst_10.BIT_WIDTH = 9;
defparam promx9_inst_10.RESET_MODE = "SYNC";
defparam promx9_inst_10.INIT_RAM_00 = 288'hAA24A5986B361F0F67B3E9E8D8720886CD67C3E1C8587F7F5BEFF7FBFDFEFF7FBFDFEE17;
defparam promx9_inst_10.INIT_RAM_01 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FAFD7EB75B6D95;
defparam promx9_inst_10.INIT_RAM_02 = 288'hEB6DBAD9568C2E134A84DAFDC7089D532DB6EB75BADD6EB75BADD7EBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_03 = 288'hEB75BADD6EB75BAFD6EB75BADD6EBF5FADD6EB75FADD6EB75FADD6EB75FAFD6EB75FADD6;
defparam promx9_inst_10.INIT_RAM_04 = 288'hEB75BADD6EB75BADD6EB75B6DD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB75BADD6;
defparam promx9_inst_10.INIT_RAM_05 = 288'hCAE572B95BADD6EB75BADD6EB55AA0A2592B3130F5DA6A240DE7149A5572BB6DB6DB6DB6;
defparam promx9_inst_10.INIT_RAM_06 = 288'hEB75B6DB6DB6DBADB6DB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6CB65B2D96;
defparam promx9_inst_10.INIT_RAM_07 = 288'hFBFDFEFF7DB6DB6DB6DB75B6DB6DB75BADD6EB75BADD6EB75BADD6DB6DBADB6EB6DB6DB6;
defparam promx9_inst_10.INIT_RAM_08 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FB85FEFF7FBFDFEE17FB85FEFF7FBFDC31F7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_09 = 288'hEBF5FADB6CAD51652CC359B0F8741E1C8366C3E9F4F678218B0F87C38C3EFD7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_0A = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_0B = 288'h68F36152995425D34BF71416333AA6576DB6EB75BAFD7FBF5FAFD7FBF5FAFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_0C = 288'hDB75BADD6EB75BADD6EB75FADD6EB75BADD6EB75BADD6EB75B6DB6EB75B6DB6DB65B2D34;
defparam promx9_inst_10.INIT_RAM_0D = 288'hDB6DB6DD6DB75BADD6EB75BADD6EB6DBADB6A9994C6633198CC644226AF29B6DB6DBADB6;
defparam promx9_inst_10.INIT_RAM_0E = 288'hDB6DB6D96CB6572B95CAE56EB75BADD6A8F35171BDF4571EBA98C2B2C90E2D39A5572B96;
defparam promx9_inst_10.INIT_RAM_0F = 288'hEB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6EB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_10.INIT_RAM_10 = 288'hFBFDFEFF7FBFDFEFF7DB6DB6DB6DB6DB6DB6DB75BADD6DB75BADD6DB75B6DD6DB6DB6DB6;
defparam promx9_inst_10.INIT_RAM_11 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDC2FF70BFDC2FF7;
defparam promx9_inst_10.INIT_RAM_12 = 288'hFBFDFEFF7FBFDFEFF7DB656A8B29669ECF87D3E1F0F66C459C8041B3E1ECF873161C63F7;
defparam promx9_inst_10.INIT_RAM_13 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_14 = 288'h94B21D3CE282CA6754BADD72BB5DB75B6DD6EB75FAFD7FBF5FEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_15 = 288'h63ED76DB6DB6DBADD6EB75BADD6EB75BADD6EB75BADD6EB6DBADB6EB6DB6DD7BB1C1D34A;
defparam promx9_inst_10.INIT_RAM_16 = 288'h9A5D72B96DB6DB6DB6EB75BADD6EB75BADD6EB75B2DAB4198CC6633198CC6633198CC643;
defparam promx9_inst_10.INIT_RAM_17 = 288'hDB6DB6DB6DB6DB6DB6CB65B2D96CAE56EB75BAD566891616B95482A60C2072440C0C1EB2;
defparam promx9_inst_10.INIT_RAM_18 = 288'hEB75B6DB6DB6DBADB6DB6DB6DB6EB6DB6DD6DB6DBADD6EB6DB2DB6CAEDBADB6DB6DB6DB6;
defparam promx9_inst_10.INIT_RAM_19 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7DB6DB6DB6DB75BADD6DB75BADD6EB75B6DB6EB75B6DB6;
defparam promx9_inst_10.INIT_RAM_1A = 288'hB3D9F0E71EBFDFF1F7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_1B = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7EBF5B6D5469D334F86C3E1E4B8720C9B0F67C3D9DC862;
defparam promx9_inst_10.INIT_RAM_1C = 288'hFBF5FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_1D = 288'h747B9E795DB6DB6DD6EB75BADD6EB75BADD6EB75FAFD7EBF5BAFD7EBF5FAFD6EBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_1E = 288'h3198CC66331A0E51B6DBF5B6DB6DB75BADD6EB75BADD6EB75BADB6DBEDBADB6CB0BD932A;
defparam promx9_inst_10.INIT_RAM_1F = 288'h045301EF39A5D72B96DB6DB6DB6DB6DBADD6EB75BADB7DB6DAE6833198CC6633198CC663;
defparam promx9_inst_10.INIT_RAM_20 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2D96CAE56EB75AA4D25861E76BD0449D6D970B65;
defparam promx9_inst_10.INIT_RAM_21 = 288'hEB75BADD6DB75B6DD6DB6DB6DB6DB6DB6DD6EB6DBADB6EB6DBADD6EB75BADB6DB6DB2DB6;
defparam promx9_inst_10.INIT_RAM_22 = 288'hFBFDC2FF7FBFDC2FF7FBFDFEFF7FBFDFEFF7DB6DB6DB6DB65B6DD6DB6DBADD6EB75B6DB6;
defparam promx9_inst_10.INIT_RAM_23 = 288'h109868D87B361D8987497DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_24 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FAFB6BAB4E5987C3E1F0FA7B3E1F4F87;
defparam promx9_inst_10.INIT_RAM_25 = 288'hEBFDFAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAFF7EBF5BAFB6DB6DBADD7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_26 = 288'h74EB56575EB6DBADD6EB75FAFD7EBF5FAFD7EBF5FADD7EBF5FAFD7EBF5FAFD7EBF5FEFD7;
defparam promx9_inst_10.INIT_RAM_27 = 288'h3198CC6633198CC6633198D07ABDBF5B6DB6DB75BADD6EB75BADD6EB6DB6DB6DB5D1D32A;
defparam promx9_inst_10.INIT_RAM_28 = 288'h65D9504A285EB92514AAE572DB6DB6DB6DB6EB6DBADD6EB75BADB7DB6D98E633198CC663;
defparam promx9_inst_10.INIT_RAM_29 = 288'hDB6DB6DB6DB75B6DD6DB6DB6DB6DB6DB6DB6DB6DB6D96CAE56EB55AA4CE8849C6B8FCE51;
defparam promx9_inst_10.INIT_RAM_2A = 288'hEB75BADD6EB75BADB6DB6DBADB6DB6DB6DB6DB6DB6DB6DB75B6DB6DB75B6DD6EB6DB6DD6;
defparam promx9_inst_10.INIT_RAM_2B = 288'hFBFDFEFF7FBFDC2FF70BFDFEFF7FBFDFEFF7FBFDFEFF7DB6DB6DB6DB6DBADD6DB75BADB6;
defparam promx9_inst_10.INIT_RAM_2C = 288'hC3E9C4105C3C970D677210B0D66B3A4FADF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_2D = 288'h9A75FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAFD6EB555A72CC3D9B4F87;
defparam promx9_inst_10.INIT_RAM_2E = 288'hEB6DBADB6EB75BADD6EB75BADD6EBF5FAFD7EBF5BADD6EB6DB6D75496B955E79230986C3;
defparam promx9_inst_10.INIT_RAM_2F = 288'hA55301ED2BAE576DB6EBEDBADB6EB75FAFD7EBF5FAFD7EBF5FADD6EBF5FAFD7EBF5FADD6;
defparam promx9_inst_10.INIT_RAM_30 = 288'h3198CC6633198CC6633198CC6633198CC6A5DB75BADD6DB6DB6DB6EB6DB6DB6DB65A66C8;
defparam promx9_inst_10.INIT_RAM_31 = 288'hE3C975C28A2BAD8669B6941E754BAE572DB6DB6DB6DB6EB6DBADD6EB75BADB6DB6550883;
defparam promx9_inst_10.INIT_RAM_32 = 288'hEB75BADD6EB6DB6DB6DB6DB6DD6DB6DB6DB6DB6DB6DB6DB6DB6D96CADD6EB559A44D87A6;
defparam promx9_inst_10.INIT_RAM_33 = 288'hEB75B6DB6EB6DB6DB6DB75B6DD6EB75BADD6EB75BADB6DB6DB6DB6DB6DB6DD6DB75B6DD6;
defparam promx9_inst_10.INIT_RAM_34 = 288'hFBFDFEFF7FB85FEFF7FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFAFF7DB6DB6DB6DB6DBADB6;
defparam promx9_inst_10.INIT_RAM_35 = 288'h9669F0F87A2D9F0F67C3E1C8242B361ECD87B359DA7F6FBFDFEFF70BFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_36 = 288'h6128A09E7AAF5BEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EB6DAEAD2;
defparam promx9_inst_10.INIT_RAM_37 = 288'hBAC53DE2871A8984C25128944C26130944A25128944A261A8D86C361B0DC6C26138D86C3;
defparam promx9_inst_10.INIT_RAM_38 = 288'h74C26960F695532BB6DB6DBADD6EB75BADD6EB75BADD6EB75BADD6EB75BADB6DB6DB6D96;
defparam promx9_inst_10.INIT_RAM_39 = 288'hDB65548633198CC6633198CC6633198CC6633198CC6E7CB6DB6DD6EB6DBADB6DB6DB2D95;
defparam promx9_inst_10.INIT_RAM_3A = 288'h9A6B986C3619234D856128B0D6C07B4A6955BAE572DB6DB6DB6DB6DB75BADD6EB6DBADD6;
defparam promx9_inst_10.INIT_RAM_3B = 288'hEB6DB6DD6DB75BADD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D96CADD6AB54;
defparam promx9_inst_10.INIT_RAM_3C = 288'hDB6DB6DB6DB6DBADD6DB75BADD6EB75B6DB6DB75BADB6EB75BADB6DB6DBADB6DB75B6DD6;
defparam promx9_inst_10.INIT_RAM_3D = 288'hFBFDFEFF7FBFDFEFF70BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAFF7DB6DB6DB6;
defparam promx9_inst_10.INIT_RAM_3E = 288'hFBF5BAD9579CB34D87C3E1F0F87103934E21B359ACCC3B3D9B0EB3EBFDFEFF7FBFDFEFF7;
defparam promx9_inst_10.INIT_RAM_3F = 288'hA642F1BEF181C5E775DB75FEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;

pROMX9 promx9_inst_11 (
    .DO({promx9_inst_11_dout_w[26:0],promx9_inst_11_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_23),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_11.READ_MODE = 1'b1;
defparam promx9_inst_11.BIT_WIDTH = 9;
defparam promx9_inst_11.RESET_MODE = "SYNC";
defparam promx9_inst_11.INIT_RAM_00 = 288'h61A8944A2821229BCE079C5A4D279BCDE6F379BCDA4B2489C4E27128140A0B2389C52250;
defparam promx9_inst_11.INIT_RAM_01 = 288'hCA8BDD30A17AC66975CB6DB6DB6DB75B6DB6EB75BADD6EB75BADD6EB75B6DB6DB65A692C;
defparam promx9_inst_11.INIT_RAM_02 = 288'hEB6DB6DD6DB65508633198CC6633198CC6633198CC6633198CC912CB75B6DB6DB6DB6DB6;
defparam promx9_inst_11.INIT_RAM_03 = 288'hCADD6AB54898235F8681C930AA251492980F59452A975CAE5B2DB6DB6DB6DB6EB75BADD6;
defparam promx9_inst_11.INIT_RAM_04 = 288'hEB75B6DD6DB6DBADD6EB75BADD6DB6DBADB6EB75BADB6DB6DB6DB6DB6DB6DB6DB6DB2D95;
defparam promx9_inst_11.INIT_RAM_05 = 288'hDAEDB6DB6DB75BADB6DB6DBADB6DB75BADD6DB6DBADD6EB75BADD6EB75BADB6EB75BADD6;
defparam promx9_inst_11.INIT_RAM_06 = 288'hFBFDFEFF7FBFDFEFF7FB85C2FF7FB85FEFF7FBFDFEFF70BFDC2FF7FBFDFEFF70BFDFEFF7;
defparam promx9_inst_11.INIT_RAM_07 = 288'hFBFDFEFF7FBFDFEFD6CABCE5986B3E1D0547D3E1ECF667220A8D66B3D9B0D8769F5BEFF7;
defparam promx9_inst_11.INIT_RAM_08 = 288'h89AC562F279A44E0D2694D2EA9148EDBEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_09 = 288'h51A8BD16D07A45A734AADD72BB6DB6DB6DB6DB75BADD6EB6DBADB6CADD4E2D279245A313;
defparam promx9_inst_11.INIT_RAM_0A = 288'hDB6DAEAC984FB8A0F3AA6576DB6DB75BADB6EB6DBADD6EB75BADD6EB6DB6DB6DB656ABE7;
defparam promx9_inst_11.INIT_RAM_0B = 288'hEB6DBADB6EB75BADB6DB6D8DC823198CC6633198CC6633198CC6633120ED5B6DB6DB6DB6;
defparam promx9_inst_11.INIT_RAM_0C = 288'hDB6DB2D95CADD6A913B2B9249041471944E3555B460D28A552EB75CB65B6DB6DB6DB6DB6;
defparam promx9_inst_11.INIT_RAM_0D = 288'hEB6DB6DD6DB75BADD6EB6DBADB6EB75BADD6DB75BADD6DB6DBADB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_11.INIT_RAM_0E = 288'hFBFDFEFF7DB6DB6DB6DB75B6DD6DB6DBADB6EB75FAFB6EB75BADD6DB6DB6DD6EB6DB6DB6;
defparam promx9_inst_11.INIT_RAM_0F = 288'hC3B4FADF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_10 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7EB655E72CC3E1F0F67C359D04E5C39020B66A3496CD46;
defparam promx9_inst_11.INIT_RAM_11 = 288'hA9BC9A2F289B49A4F289BC9E51399B49E51399BCF6D95DAFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_12 = 288'hE3A8ACBAE38BCEEB75CAEDB6DB6DB75BADD6EB75BADD6EBF5FAFD6EB6DB6CF358BCDA513;
defparam promx9_inst_11.INIT_RAM_13 = 288'hDB6DB6D96CAB22123048C4EA975DB6DB6DB6EB75BADB6EB6DBADB6DB6DBADB6DB65B2B35;
defparam promx9_inst_11.INIT_RAM_14 = 288'hDB6DB6DB6DB6DBADB6EB75BADB6EB6DAA8633198CC6633198CC6633198CC66331C232DB6;
defparam promx9_inst_11.INIT_RAM_15 = 288'hDB6DB6DB6DB6DB2D95BADD66889925960924E320A88EAD7145A513AA5D72B95CB6DB6DB6;
defparam promx9_inst_11.INIT_RAM_16 = 288'hEB75BADB6DB6DBADD6EB75BADD6DB6DBADD6EB75BADD6DB75BADD6EB6DBADD6EB75B6DB6;
defparam promx9_inst_11.INIT_RAM_17 = 288'hFBFDFEFF7FBFDFEFF7DB6DB6D96DB75BADD6EB75BADD6EB75BADB6DB6DB6DD6EB75BADB6;
defparam promx9_inst_11.INIT_RAM_18 = 288'hB318A8D66B359D65D6EB7DFEE17FBFDFEFF7FBFDFEE17FB85FEFF7FBFDFEFF8FC7DFEE17;
defparam promx9_inst_11.INIT_RAM_19 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5B2B1385E9ECF873149ACD46B359B0F05;
defparam promx9_inst_11.INIT_RAM_1A = 288'h9A44DA4F289C4920D168839A2F2892C5A4F289B49A4F389C4E27339A3CFADF7FBFDFEE17;
defparam promx9_inst_11.INIT_RAM_1B = 288'hBAF3D44E3C724A6975CAEDB6DB6DB75BADD6EB75BADD7EB75FADD7EBF5FADD6EB6D9E4F3;
defparam promx9_inst_11.INIT_RAM_1C = 288'hC66DB6DD6CB6D6EB09741C52514BAE5B2DB6DB6DB6DD6EB75BADB6DB6DB6DD6DB6DB6D96;
defparam promx9_inst_11.INIT_RAM_1D = 288'hCB6DB6DB6DB6DB6DD6DB6DBADD6EB75BADD6EB6DB2D8A41A0CC6633198CC6633198CC483;
defparam promx9_inst_11.INIT_RAM_1E = 288'hDB6DBADB6DB6DB6DB6DB65B2D75BAD501EC371E1B0B6551E9A17CE38B4E2954BAE572B96;
defparam promx9_inst_11.INIT_RAM_1F = 288'hEB75BADB6DB75BADB6EB75BADD6DB75B6DB6EB75B6DB6EB75BADD6DB75BADD6EB6DBADB6;
defparam promx9_inst_11.INIT_RAM_20 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7DB6DB6DB6DB6DBADB6DB6DBADD6DB75BADD6DB75BADB6;
defparam promx9_inst_11.INIT_RAM_21 = 288'hB351B0E414151A8D66B328F0ED2EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_22 = 288'h89D53EE17FBFDC2FF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFAD9589C330D66C3D1B0D86;
defparam promx9_inst_11.INIT_RAM_23 = 288'hDB4D1E51379C4D62B17944A6733AA551E4B1693C920F27924162F2892462734BA4CE2713;
defparam promx9_inst_11.INIT_RAM_24 = 288'hCB5D66924511A46134BAE5B2DB6DB6DB6DD6EB75BADD6EB75BADD7EB75FADD7EBF5FADD6;
defparam promx9_inst_11.INIT_RAM_25 = 288'h3198CC8D1CB6DB6DB6BB52E547148C52AB96DB6DB6DB6DB6DB6DD6EB75BADB6DB6DB6DB6;
defparam promx9_inst_11.INIT_RAM_26 = 288'hBAE572DB6DB6DB6DB6DB6DB6DB6DB75BADD6EB75B6DD6EB6DB2D745218CC6633198CC663;
defparam promx9_inst_11.INIT_RAM_27 = 288'hEB75BADB6EB6DB6DB6DB6DB6DB6CB65AEB75BAACA06A35128A06A261C2F5C5079CD2AB75;
defparam promx9_inst_11.INIT_RAM_28 = 288'hEB75BADD6DB6DB6DD6DB75B6DD6DB75B6DB6DB75B6DD6EB75BADD6EB75BADD6EB6DBADD6;
defparam promx9_inst_11.INIT_RAM_29 = 288'hFBFDFEE17FBFDFEFF7FBFDFEFF7FBFDFEFD7DB6DB6DB6DB75F6DD6EB75BADD6EB75BADB6;
defparam promx9_inst_11.INIT_RAM_2A = 288'hC3D9A0B258290ACD86B3D9ACC417251ACD475975BEDF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_2B = 288'h89BC9E533AA3CFADF7FBFDC2FF70BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF6DB44E1966;
defparam promx9_inst_11.INIT_RAM_2C = 288'hEBF5FADB69A44E27138944E6974CAEDBADD6EB75BADB6EB6DB6B95CAE56E93379245E513;
defparam promx9_inst_11.INIT_RAM_2D = 288'hDB6DB2D75D730D87AE695D72BB6DB6DB6DD6EB75BADD6EB75BADD6EB75BADD7EBF5BAFD7;
defparam promx9_inst_11.INIT_RAM_2E = 288'h3198CC66331B16EB96DB6DB2CF38494162F3AAE572DB6DB6DBADB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_11.INIT_RAM_2F = 288'h8A552EB75CB65B6DB6DB6DB6DB6DB6DB6DB6DB75BADD6DB75B6DB6DB6DB6D9626A0CC663;
defparam promx9_inst_11.INIT_RAM_30 = 288'hEB6DBADD6EB6DBADD6DB6DB6DB6DB6DB6DB6CB656EB559A49249E78241248A285EB8A0D3;
defparam promx9_inst_11.INIT_RAM_31 = 288'hEB75BADD6EB6DB6DB6EB75B6DD6EB75BADD6EB6DBADB6DB75BADD6EB75BADD6EB75BADB6;
defparam promx9_inst_11.INIT_RAM_32 = 288'hFBFDFEFF70BFDFEFF70BFDFEFF7FBFDFEFF7FBFDFEFF7DB6576DB6DB6DBADD6DB6DBADD6;
defparam promx9_inst_11.INIT_RAM_33 = 288'hEB65A26CBB359A8D66B359A8F87C31050566A359A8C41B324BEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_34 = 288'hEB656A8F248A45E4F299BC9E4D20BFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_35 = 288'hEBF5FAFD7EBF5B6D75794CEA93399E536DD6EB7DFADF7FBFDFEFF7FBFDFEFF7FBFDFADD6;
defparam promx9_inst_11.INIT_RAM_36 = 288'hDB6DB6DB6CB65A0882249C66995CB6DB6DB6DB6DBADD6EB75BADD6EB75BADD7EBF5FAFD7;
defparam promx9_inst_11.INIT_RAM_37 = 288'hDAA11066331989068489E5F6DB6CB6D550C948ACA6975CAEDB6DB6DB6DB6DB6DB75B6DB6;
defparam promx9_inst_11.INIT_RAM_38 = 288'hB68C16513AADD72B96CB6DB6DB6DB6DB6DB6DB6DB6DB6EB75B6DD6EB6DBADB6DB75BADB7;
defparam promx9_inst_11.INIT_RAM_39 = 288'hEB75B6DD6EB75BADB6DB6DB6DB6DB6DB6DB6DB6DB6DB6CADD6EB54A2B0E494571E154428;
defparam promx9_inst_11.INIT_RAM_3A = 288'hEB75BADD6EB75BADD6EB75BADB6DB75BADB6EB6DBADB6EB75BADB6EB75BADD6EB75BADD6;
defparam promx9_inst_11.INIT_RAM_3B = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FB85FEFF7FBFDFEFF7FBFDFEFF7CB6DB6DB6DB6DB6DD6;
defparam promx9_inst_11.INIT_RAM_3C = 288'hFBFDFEFF7FBF5B6D3475D9B0D66C3D99C800A359ACD66A28850745A351863D6FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_3D = 288'hFBFDFEFF7FBF5BADD6DAC4D62F268BCA2733697DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_3E = 288'hEBF5FAFD7EBF5FAFD6DB6DB2CF389C4E2713CAF5BADF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_11.INIT_RAM_3F = 288'hDB6DB6DB6DB6DAEA9261A071AF3BAE5B6DB6DB6DB6DB6EB6DBADD6EB75BADD6EB75BADD6;

pROMX9 promx9_inst_12 (
    .DO({promx9_inst_12_dout_w[26:0],promx9_inst_12_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_25),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_12.READ_MODE = 1'b1;
defparam promx9_inst_12.BIT_WIDTH = 9;
defparam promx9_inst_12.RESET_MODE = "SYNC";
defparam promx9_inst_12.INIT_RAM_00 = 288'hDB6DB6DB6DB6548A834229E2596DB6DB2DB6694A5A4B189D532B96DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_01 = 288'hA230A092CF7ACA2754BADD72B96DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DBADB6EB75BADB6;
defparam promx9_inst_12.INIT_RAM_02 = 288'hEB75BADD6EB75BADD6EB75BADD6DB6DB6DB6EB6DB6DB6DB6DB2D96BADD6686992021C6C3;
defparam promx9_inst_12.INIT_RAM_03 = 288'hDB6DBADD6EB75BADD6EB75B6DD7EB6DB6DB6EB75B6DD6DB75BADD6EB75BADB6DB75BADB6;
defparam promx9_inst_12.INIT_RAM_04 = 288'hFB75BEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_05 = 288'hFBFDFEFF7FBFDFEFF7FBFDFADB68A3AE8D66B35168D66B351B0C2020D1A8D2582A8E8FEF;
defparam promx9_inst_12.INIT_RAM_06 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7EBEDB2B1258BC9E53389CD1E795FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_07 = 288'hEB75BADD6EB75FAFD7EBF5BADD6DB5D5E734BA44DE554DB75BAFD7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_08 = 288'hEB6DB6DB6DB6DB6D96BAB2D8585184D2EBB6DB6DB6DB6DB75BADD6EB75B6DD6EB75BADD6;
defparam promx9_inst_12.INIT_RAM_09 = 288'hDB75B6DD6DB6DB6DB6DB6DB6D74BA6DB2DB6DB6DAAB8C84AC9A534BAE5B6DB6DB6DB6DD6;
defparam promx9_inst_12.INIT_RAM_0A = 288'h51289470381A8A17CE38BCE6955BAE572B96DB6DB6DB6DB6DB6DB6DB6DB6DB6EB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_0B = 288'hEB6DBADB6EB75BADD6EB6DBADD6EB75B6DD6EB6DB6DB6DB6DB6DB6DB65B2D95BAD579EA2;
defparam promx9_inst_12.INIT_RAM_0C = 288'hDB6DB6DB6DB6DBADD6DB75BADD6EB75BADD6EB75BADB6EB6DBADD6DB6DBADD6EB75BADD6;
defparam promx9_inst_12.INIT_RAM_0D = 288'h4151ACD66C775BAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF70BFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_0E = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFD6DB5519766B359A8D66829824BA730C164AC3;
defparam promx9_inst_12.INIT_RAM_0F = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FAD95793C9E4F27944EA933CAFDFEFF7;
defparam promx9_inst_12.INIT_RAM_10 = 288'hEB75BADD6EB75BAFD6EB75BADD6EB75B6DB6DB4D2271399C4EE9B6EB75FAFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_11 = 288'hDB6DB6DB6DB6DB6DB6DB65AEA08511A56555BAE5B6DB6DB6DB6DB6DB75BADB6EB75BADD6;
defparam promx9_inst_12.INIT_RAM_12 = 288'hDB6DB6DB6DB6DB6DB6DB75B6DB6DB6DB6DB6DB6DB6DB6CB5D7192B58BCEA975CB65B6DB6;
defparam promx9_inst_12.INIT_RAM_13 = 288'hAAAC9876571A8945A551AAB1A50694D2AB75CAE5B2D96DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_14 = 288'hDB75B6DD6EB75B6DD6EB75BADD6EB75BADD6EB6DB6DB6DB6DB6DB6DB6DB6D96CB65B2B75;
defparam promx9_inst_12.INIT_RAM_15 = 288'hFBFDFEFF7DB6DB6DB6DB6DB6DB6EB75B6DD6DB75B6DD6EB6DBADB6EB6DBADD6DB6DBADD6;
defparam promx9_inst_12.INIT_RAM_16 = 288'hA2988C525A351A8D66A3433AFD6FBFDFEFF7FBFDFEFF7FBFDC2FF7FBFDFEE17FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_17 = 288'hCAFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7EBEDAA8CBA35168C009359A4D45;
defparam promx9_inst_12.INIT_RAM_18 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFD7DB5D2269089449E533;
defparam promx9_inst_12.INIT_RAM_19 = 288'hEB75B6DD6EB75BADD7EBF5BADD6EB75BADD6EB75BADB6CAD5227139A4CF2BD6FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_1A = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6BAF1D450B89DD76DB6DB6DB6DB6DB6DB6DB6EB75BADD6;
defparam promx9_inst_12.INIT_RAM_1B = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DD6DB6DB6DB6DB6DB6DB6DB6DB2D96CA9C2969179D52EB96;
defparam promx9_inst_12.INIT_RAM_1C = 288'hCB656EB559A392090461D1090A2D2D33DEB289D56EB75BAE5B6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_1D = 288'hEB6DB6DD6DB6DB6DD6EB75BADD6EB75B6DB6EB75BAFD6EB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_1E = 288'hFBFDFEFF7FBFDFADF7DB6DB6DB6DB6DBAFD6EB75BADD6EB75F6DB6EB75B6DD6EB75B6DB6;
defparam promx9_inst_12.INIT_RAM_1F = 288'hA2C968A62928A04104935994746A351A19B6EBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_20 = 288'h483CA273389E57EFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5B6D54555168D45;
defparam promx9_inst_12.INIT_RAM_21 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5BAD33;
defparam promx9_inst_12.INIT_RAM_22 = 288'hEB75BADD6EB6DBADD6DB75FADD6EB75BADD6EB75FADD6EB75BADB6CAD522754AA3CF6BD6;
defparam promx9_inst_12.INIT_RAM_23 = 288'hAADD72DB6DB6DB6DB6DB6DB6DB6DB6DB2DEF6132A2975CB6DB6DB6EB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_24 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6DB6DB6DB6DB6DB6DB6DB6DB2D959A5AD22F3;
defparam promx9_inst_12.INIT_RAM_25 = 288'hDB6DB6D96CADD6EB3471F1F8EC381C9102C285F3D22F39A556EB95CAE5B6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_26 = 288'hEB75BADB6DB6DB6DD6DB6DB6DD6EB75BADB6EB75B6DB6EB75BADB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_27 = 288'hFB85C2FF7FBFDFEFF7FBFDFEFF7DB6DB6DB6DB6DBAFD6DB6DBADD6DB75BADD6EB6DB6DD6;
defparam promx9_inst_12.INIT_RAM_28 = 288'h9A2AA4B45930024CE4A351A8D46725194746A351A8CABEB75BEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_29 = 288'hFBF5FAF9599B462734AA3CFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5BADB6;
defparam promx9_inst_12.INIT_RAM_2A = 288'h99CCF6BD6EB75FAFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_2B = 288'hEB6DB6DB6DB6DB6DD6EB75BADB6EB75BADD6EB75BADD6EB75BADD6EB75B6DB6CAC4E2713;
defparam promx9_inst_12.INIT_RAM_2C = 288'h849C1A574BAE5B6DB6DB6DB6DB6DB6DB6DB6CB4D187048A6572DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_2D = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6CB65AEB55;
defparam promx9_inst_12.INIT_RAM_2E = 288'hDB6DB6DB6DB65B2D95BADD6ABE76149146C3A2C0D44EAC7141A534AADD72B96CB65B6DB6;
defparam promx9_inst_12.INIT_RAM_2F = 288'hEB75B6DB6DB75BADB6DB75B6DB6DB6DBADB6DB75BADB6EB75B6DD6EB75BADB6DB75B6DB6;
defparam promx9_inst_12.INIT_RAM_30 = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBF5FAFD7DB6DB6DB6DB6DB6DD6EB75BADD6EB75BADB6;
defparam promx9_inst_12.INIT_RAM_31 = 288'hFBF5BADD6DB5555525A35168D469349A4DC740A0E8D66A3518C54614F5BAFD7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_32 = 288'hFBFDFEFF7FBF5BADD6BAAC626F289C4FADF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_33 = 288'hCAC4DA51379D532BD6EBF5FAFD7EBF5FEFF7FBFDFAFD7FBFDFAFD7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_34 = 288'hDB6DB6DB6DB6DB6DB6EB6DB6DD6EB75B6DD6EB75BADD6EB75BADD6EB75BADD7EB75B6DB6;
defparam promx9_inst_12.INIT_RAM_35 = 288'hDB5D72AE938C4EAB75CB6DB6DB6DB6DB6DB6DB6DB6D9589A8B1B75CB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_36 = 288'hDB65B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_37 = 288'hDB6DB6DB6DB6DB6DB6CB65B2B75BAD52DAA392B8D86C3F3A88916C07A462754BADD72B96;
defparam promx9_inst_12.INIT_RAM_38 = 288'hEB75BADD6DB6DB6DB6DB75BADB6DB6DB6DB6DB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_39 = 288'hEB7DFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFADD6DB6DB6DB6DB6DB6DB6DB75BADD6;
defparam promx9_inst_12.INIT_RAM_3A = 288'hFBFDFEFF7FBF5FADD6EB6DAAAAA92D1A8CE4A2B0C8325B35168B465190A4D45928A76DF7;
defparam promx9_inst_12.INIT_RAM_3B = 288'hFBFDFEFF7FBFDFEFF7FBFDFAFD6DB54CE0B17944E26F2FBFDFEFF7FBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_3C = 288'hDB6DB6D95BAB4A273489D53ADD6EBF5FAFD7FBF5FEFF7FBFDFAFD7EBFDFEFF7FBFDFEFF7;
defparam promx9_inst_12.INIT_RAM_3D = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6EB75BADD6EB6DBADD6EB75BADD6EB75BADD6;
defparam promx9_inst_12.INIT_RAM_3E = 288'hDB6DB6D96CADD50E0F58CD2EB96CB6DB6DB6DB6DB6DB6DB65AEA91517BEEBB6DB6DB6DB6;
defparam promx9_inst_12.INIT_RAM_3F = 288'hBAE572B96DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;

pROMX9 promx9_inst_13 (
    .DO({promx9_inst_13_dout_w[26:0],promx9_inst_13_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_27),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_13.READ_MODE = 1'b1;
defparam promx9_inst_13.BIT_WIDTH = 9;
defparam promx9_inst_13.RESET_MODE = "SYNC";
defparam promx9_inst_13.INIT_RAM_00 = 288'hDB6DB6DB6EB6DB6DB6DB6DB6DB6CB6572B75AAA4544C361B0E8A6950D1257CE48BCE6955;
defparam promx9_inst_13.INIT_RAM_01 = 288'hEB6DBADB6DB6DB6DB6DB6DB6DD6EB6DB6DB6DB75BADB6EB6DB6DB6DB6DB6DB6DB6DBADD6;
defparam promx9_inst_13.INIT_RAM_02 = 288'h314978FB6EBFDFEFF7FBFDFEFF7FBFDFEE17FBFDFEFF7FBF5BEFD6CB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_03 = 288'hFBFDFEFF7FBFDFEFF7EB75BADD6EB75F6D5475C168D46A351A8B46A2D990241935164B46;
defparam promx9_inst_13.INIT_RAM_04 = 288'hEBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFD6EB65626D17944EA933CAFDFEFF7FBFDFEFF7;
defparam promx9_inst_13.INIT_RAM_05 = 288'hEB75BADD6DB6DB6D9589BC9E4F2794D36DD6EBF5FAFD7EBFDFEFD7EBF5FEFF7FBF5FEFD7;
defparam promx9_inst_13.INIT_RAM_06 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6DB6DB6DD6EB75BADD6;
defparam promx9_inst_13.INIT_RAM_07 = 288'hDB6DB6DB6DB6DB6D95BABA696919A5D72B96DB65B6DB6DB6DB6DB6DB5D564C307D532DB6;
defparam promx9_inst_13.INIT_RAM_08 = 288'h69452A975BAE572D96DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_09 = 288'hDB6DBADD6DB6DB6DB6DB6DB6DB6DB6DB2D96CADD6EB7579B098745C3516CAC25132F5C50;
defparam promx9_inst_13.INIT_RAM_0A = 288'hDB6DB6DD6EB75BADD6EB6DB6DB6DB6DB6DB6DB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_0B = 288'hA351A4A40A2D164D86DB75BEFF7FBFDFEFF7FBFDFEFF7FBFDFEFD7FBF5FEFD7CB65B6DB6;
defparam promx9_inst_13.INIT_RAM_0C = 288'hFBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFADD6EB75BEDD6BAAAE4B46A35168D2520496CD25;
defparam promx9_inst_13.INIT_RAM_0D = 288'hEBF5FAFF7EBFDFEFF7FBFDFEFD6FB7DFEFF7FBFDFADF7EB6DAA89079349E4F2DAF5BEFF7;
defparam promx9_inst_13.INIT_RAM_0E = 288'hEB75BADD6EB75B6DD6DB6DB6D9589AC5A4F289C4F6BD6EB75FAFD7EBF5FEFF7FBF5FAFD7;
defparam promx9_inst_13.INIT_RAM_0F = 288'h9A5D76DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6EB6DB6DB6DB75B6DB6DB75BADD6;
defparam promx9_inst_13.INIT_RAM_10 = 288'hDB6DB6DB6DB6DB6DB6DB65B2B7517CA8E314BAE572DB6DB6DB6DB6DB6DB6D96BABCD45EF;
defparam promx9_inst_13.INIT_RAM_11 = 288'h44DB45EB289CD2EB75CAE5B2DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_12 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB65B2D95BAD56AB34E340E06C38241248A2;
defparam promx9_inst_13.INIT_RAM_13 = 288'hCAE576DB6DB6DB6DB6DB75B6DB6DB6DB6DB6DB6DB6DB6EB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_14 = 288'hA2D168D66109060B46A34968B05B3657AFD7EB75FEFF7FBFDFEFF7FBFDFAFF7FBF5FAFD6;
defparam promx9_inst_13.INIT_RAM_15 = 288'h79553EFF7FBFDFEFF7FBFDFEFF7FBFDFADD6EB7DFADF7EB7DFADD6DB5555725A2D190725;
defparam promx9_inst_13.INIT_RAM_16 = 288'hEBF5FAFD7EBF5FAFD7EBFDFEFF7FBFDFADF7FBFDFEFF7EB7DFEFD6EB75B2B1338241E513;
defparam promx9_inst_13.INIT_RAM_17 = 288'hDB6DB6DB6EB75BADD6DB6DB6DB6DB6DB6DB6BAC4DE51299CD1E5B6EB75FAFD7EBF5FAFD7;
defparam promx9_inst_13.INIT_RAM_18 = 288'h9A28B9F13BAE5B2DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_19 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6CB65AEB34849C1E775BAE5B2DB6DB6DB6DB6CB65B2B75;
defparam promx9_inst_13.INIT_RAM_1A = 288'h71F9D45A6A67B922F39A556EB75CAE5B2DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_1B = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D96CB65B2B75BAD56290471B8D4586;
defparam promx9_inst_13.INIT_RAM_1C = 288'hEB75FAFD6CB6576DB6DB6DBADB6DB75B6DD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_1D = 288'h92D168B469351442E4C31860925A318A4D45A2D9F6DD6FB75FEFF7FBFDFEFF7FBFDFEFD7;
defparam promx9_inst_13.INIT_RAM_1E = 288'h793C5E533AA44FADF7FBF5BEFF7FBFDFEFF7FBF5BADD6EB75BADF7EB75BEFD6EB6DAEAEB;
defparam promx9_inst_13.INIT_RAM_1F = 288'hEBF5FAFD7EBF5FAFD7EBFDFAFD7FBF5FAFF7FBFDFADF7EB75BEFF7EB7DFEFD6EB75B6D75;
defparam promx9_inst_13.INIT_RAM_20 = 288'hDB6DB6DB6DB6DB6DB6EB75BADB6EB6DB6DB6DB6DBADB6CAD51E4F279CCDE795EB75FAFD7;
defparam promx9_inst_13.INIT_RAM_21 = 288'hCB656EB3451535A755CAE5B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_22 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB65B2D96CB65669093834AEB95CB65B6DB6DB6DB2DB6;
defparam promx9_inst_13.INIT_RAM_23 = 288'hF3B8D45441428986EBD7141A514AA556EB95CAE5B2DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_24 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D96CADD6EB55AA4D092C3;
defparam promx9_inst_13.INIT_RAM_25 = 288'hFBFDFAFF7FBF5FADD6CB6DB2DB6DB6DB6DB6DB6DB6DB6EB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_26 = 288'hEB75BAD54864168B46104168D2592D16CCA292D160B25A351B0D76FB7DFADF7EB7DFEFF7;
defparam promx9_inst_13.INIT_RAM_27 = 288'hEB75FADB689B45A2F2893CBADD6EB75BADF7EB7DFEFF7FBF5BEFF7EB75BADD6EB75BADD6;
defparam promx9_inst_13.INIT_RAM_28 = 288'hEB75BADD7EBF5FAFD7EBF5FAFD7EBF5FAFD7FBF5FAFD7EBF5FADD6EB7DFEFD6EB7DFADD6;
defparam promx9_inst_13.INIT_RAM_29 = 288'hDB6DB6DB6DB6DB6DB6DB75B6DD6EB75BADB6DB6DBADD6DB6DB6DB6DAD51A4D269349E734;
defparam promx9_inst_13.INIT_RAM_2A = 288'hCB65B2D95CADD6A9E7B2A4A6975CAE5B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_2B = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2D96BAD5191CE59552AB96CB65B6DB6;
defparam promx9_inst_13.INIT_RAM_2C = 288'h9A7BDC6A361D130DE761A89556D182CA2734AA5D6EB95CAE5B6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_2D = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB65B2B75BAD56A954;
defparam promx9_inst_13.INIT_RAM_2E = 288'hFBFDFEFF7FBFDFEFF7FBF5FEFD6DB65B6DB6DB6DB6DB6DB6DB6DD6DB6DB6DB6EB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_2F = 288'hFBFDFADD6EB75BADB6BAC320B2592D168B45934164D243051A8B46A33968D87AAF5BADD6;
defparam promx9_inst_13.INIT_RAM_30 = 288'hFBF5BADD6EB75BADB6BA34920F299C4FADD6EB7DFEFF7FBF5BADD6EB75BADD6EB75BADD6;
defparam promx9_inst_13.INIT_RAM_31 = 288'h6944E6913AA6DBAFD7EBF5FAFD7FBFDFAFD7EBF5FAFF7FBFDFADD6EB75BADD6EB75BEFF7;
defparam promx9_inst_13.INIT_RAM_32 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6EB75BADB6EB6DB6DB6DB5D668F2;
defparam promx9_inst_13.INIT_RAM_33 = 288'hCB65B6DB6DB65B2D95BAD54A2C228452EB95CB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_34 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB65B2B75BAF3614719A5D72B96;
defparam promx9_inst_13.INIT_RAM_35 = 288'hAAD52691438B8D87040451649C6408A299EF48BCE6954AADD72B95CAE5B6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_36 = 288'hDB6DBADB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D96CB656EB75;
defparam promx9_inst_13.INIT_RAM_37 = 288'hB3557EFD6FBF5BEFF7FBFDFAFD7EBF5FAFD6CB65B6DB6DB6DB6DB6DB6DB6DD6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_38 = 288'hFBFDFADD6EB75BADD6EB75BADD6DB5D6192592D160B25A28824B269359B0D66105168B45;
defparam promx9_inst_13.INIT_RAM_39 = 288'hEB7DFADD6FBF5BADD6FBF5BADB6CACCE2513BA5D227D6EB75BEFD6FBFDFEFD6EBF5BEFF7;
defparam promx9_inst_13.INIT_RAM_3A = 288'hDB656A8F268BC9A513AA6DBADD6FBF5FAFD7EBF5FAFD7EBFDFADD6EB75BADD6EB75BADD6;
defparam promx9_inst_13.INIT_RAM_3B = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6DB6DBADD6EB6DB6DD6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_3C = 288'hBADD72B96CB65B6D96CB65B2D75AAC51863079D52EB95CB65B6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_3D = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D96DB6DB2B75AA424E113;
defparam promx9_inst_13.INIT_RAM_3E = 288'hAAD5269349A45226B261B8C52C351C0F8CA28242F5C5169C526954AADD72B95DB6DB6DB6;
defparam promx9_inst_13.INIT_RAM_3F = 288'hEB75B6DB6DB6DBADB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2D75;

pROMX9 promx9_inst_14 (
    .DO({promx9_inst_14_dout_w[26:0],promx9_inst_14_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_29),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_14.READ_MODE = 1'b1;
defparam promx9_inst_14.BIT_WIDTH = 9;
defparam promx9_inst_14.RESET_MODE = "SYNC";
defparam promx9_inst_14.INIT_RAM_00 = 288'hA349A8B6631599A7D6EB7DFEFF7FBFDFEFD7EBF5BADD6CB65B6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_01 = 288'hEB75BADD6EB75BADD6EB75BADD6EB75BADD6EB6DAEB0C824968D46A351ACD46A340C42E4;
defparam promx9_inst_14.INIT_RAM_02 = 288'hEB75BADD6EB75BADD6EB75BEFF7EB75BADB6CACCE2513A9D5267D6EB75BADF7FBF5BEFD6;
defparam promx9_inst_14.INIT_RAM_03 = 288'hEB75BADB6DB6DAEAF258B45A4F2793CBADD6EB75FAFF7EBF5FEFD6EB75BADD6EB7DFEFD6;
defparam promx9_inst_14.INIT_RAM_04 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6EB75B6DB6DB6DB6DB6DB75B6DD6;
defparam promx9_inst_14.INIT_RAM_05 = 288'h7413DA554CAE572B96DB65B2D96CB65AEB559A1871AB29A5572B96CB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_06 = 288'hCB65B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2DB6DB6DB2DB6DB65AEB34;
defparam promx9_inst_14.INIT_RAM_07 = 288'hCAE56A954AA44E271379B492345D340DC6A3C29A104A26563460B289CD2A955BADD72B95;
defparam promx9_inst_14.INIT_RAM_08 = 288'hDB6DBADB6DB75B6DB6DB6DB6DD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2B96;
defparam promx9_inst_14.INIT_RAM_09 = 288'h61D1A09259351840C3A35168C30EB75BADD6FBFDFEFF7EBF5BEDD6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_0A = 288'hEB75BEFD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75B6D75A64964B2592D9A4C61;
defparam promx9_inst_14.INIT_RAM_0B = 288'hFBF5BADD6EB7DFEFD6EB75BADD6EB75BADF7FBF5BADB6CAD4E251399CD32BD6EB75BADD6;
defparam promx9_inst_14.INIT_RAM_0C = 288'hDB6DB6DB6EB75BADB6DB6DB2B7489A4162F299C4DE5D6EB75BADD7FBFDFADD6EB75BADD6;
defparam promx9_inst_14.INIT_RAM_0D = 288'hDB6DB6DB6DB65B2DB6DB6DB6DB6DB65B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_0E = 288'hCB5D6EBEE952466975CAE572B96CB65B2D96CADD6EB34245952313AADD72B95CB65B6DB6;
defparam promx9_inst_14.INIT_RAM_0F = 288'hBAE572B96CB65B2DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6CB6DB6D96;
defparam promx9_inst_14.INIT_RAM_10 = 288'hCAE56EAA8532990C6532A18CC8817A470AA25130B0BA6C34914489A67BD22F38A4D2A955;
defparam promx9_inst_14.INIT_RAM_11 = 288'hDB6DB6DB6DB75B6DB6DB6DB6DD6EB75B6DB6DB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_12 = 288'hA28868B26A35164D4620A0E8D46A2D15C946B6EDBEDD6FBF5BAFD7EB75BEDD6CB5D6EB95;
defparam promx9_inst_14.INIT_RAM_13 = 288'hEB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADB6BACB20B25;
defparam promx9_inst_14.INIT_RAM_14 = 288'hEB75BADD6EB75BADD6FBF5BEDF6EB75BADD6EB75BADD6EB75B6DB5AA44DE554BA4CF6DD6;
defparam promx9_inst_14.INIT_RAM_15 = 288'hDB6DB6DB6DB75B6DB6DB75BADB6DB6DB6D96BAC4D62D1693C9E533BAF5BADD6FBF5FADD6;
defparam promx9_inst_14.INIT_RAM_16 = 288'hCB65B6D96CB6DB6DB6DB6DB6D96DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_17 = 288'hDB6DB2D95CADD669091844EE975CAE572B96CB65B2B95CADD6A8D3511C5E754BAE572D96;
defparam promx9_inst_14.INIT_RAM_18 = 288'h9A4D2A955BAE572B95CB65B2DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2DB6;
defparam promx9_inst_14.INIT_RAM_19 = 288'hDB65B6B969999D0A8542A990A6532A150A8602B0986C2A26160904F32070CEBD714164F3;
defparam promx9_inst_14.INIT_RAM_1A = 288'hDB65B6DB6DB6DB6DB6DB6DB6DD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2DB6;
defparam promx9_inst_14.INIT_RAM_1B = 288'hDB5D2992592C968B4592A8D0545B30824D4682B128D46B33AF6DD6EB75BADD6EB75BADD6;
defparam promx9_inst_14.INIT_RAM_1C = 288'hA9D53ADD6EB75BADD6EB75BADF7EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75B6DD6;
defparam promx9_inst_14.INIT_RAM_1D = 288'hEB75BADD6FBF5BEFD6EB7DFEFD6EB75BADD6EB75BADF7FBF5BADD6EB75B6D95899C22513;
defparam promx9_inst_14.INIT_RAM_1E = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DBADB6EB6DBADB6CADD1A2B168AC5A4F2793CBADD6;
defparam promx9_inst_14.INIT_RAM_1F = 288'hBAE572D96CB65B6D96DB65B6DB6DB6DB6D96DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_20 = 288'hDB65B6DB6DB6DB2B95BAD5151AD49552EB75CAE572B95CAE572D95BAD5628A3282CA6955;
defparam promx9_inst_14.INIT_RAM_21 = 288'hF79C5A6F38A4D26955BAE572B95CB65B2D96CB6DB6DB6DB6DB6D96DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_22 = 288'hDB6DB6D96CB65AEB6C32A150A8542A150A8542A150A055130DC7C78238D85E751B0D956D;
defparam promx9_inst_14.INIT_RAM_23 = 288'hEB75BADD6CB65B6DB6CB6DB6DB6DB6DB6DB6DB6DB6DB6EB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_24 = 288'hEB75BADD6EB6DA696D82C964CC451D984325A2D1A8D05A28028B4592D1853B6EB75BADD6;
defparam promx9_inst_14.INIT_RAM_25 = 288'h89C4E6733AA6D7ADD6EBF5BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6;
defparam promx9_inst_14.INIT_RAM_26 = 288'h89BCBADD6EB75BEFF7FBFDFEFD6EB7DFEFF7EB75BADF7EB75BADD6FBF5BADD6EB6DB2B33;
defparam promx9_inst_14.INIT_RAM_27 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DBADD6DB75BADB6DB6D6EB1258A4162F2;
defparam promx9_inst_14.INIT_RAM_28 = 288'h5944EAB75BAE572B96CB6DB6D96CB6DB6D96DB6DB6DB6CB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_29 = 288'hDB6DB6DB6DB6DB6D96DB6572B75BAD4E12509A5532B95CAE572B95CAE5B2D75BACD34C48;
defparam promx9_inst_14.INIT_RAM_2A = 288'hD211E57AE18245A6F38A4D2A955BADD72B95CAE5B2DB6DB6DB6DB6DB6DB6DB6CB65B6DB6;
defparam promx9_inst_14.INIT_RAM_2B = 288'hDB6DB6DB6CB65B2D96CADD5D26542A150A8542A150A8542A148AC261E9B0AC361B8C1025;
defparam promx9_inst_14.INIT_RAM_2C = 288'hDB75BADD6EBF5BADD6CAE572DB6DB6DB6DB6DB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_2D = 288'hEB75BADD6EB75BADD6EB75B6D55B6C964B4592C964B25A34974C4151C968B46928828DE8;
defparam promx9_inst_14.INIT_RAM_2E = 288'hDAE56A91289CCE6754AA75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6;
defparam promx9_inst_14.INIT_RAM_2F = 288'h999C162B168BCA26D2DAF5BAFD7EBFDFEFF7EB75BADF7FBFDFADD6FBF5BEFD7EB75BADB6;
defparam promx9_inst_14.INIT_RAM_30 = 288'hDB6DB6DB6DB6DB2DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6DB6DB6DD6DB6DB6B95;
defparam promx9_inst_14.INIT_RAM_31 = 288'hAA3CD449179CD2EB75CAE572D96DB65B2D96CB65B2DB6CB6DB2D96CB6DB2D96DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_32 = 288'hDB65B2D96DB6DB6DB6DB6DB6DB6CAE572B75AA2A3DAF3AADD72B95CAE572B95CAE56EB75;
defparam promx9_inst_14.INIT_RAM_33 = 288'hD3698CC8552A150F8C1824564D389CD26955AADD72B95CB65B2D96DB6DB6DB6DB6DB6D96;
defparam promx9_inst_14.INIT_RAM_34 = 288'hDB6DB6DB6DB6DB6DB6DB65B2D95BADAD0C8552A150A8542A150A854299A46E3D338DC6E3;
defparam promx9_inst_14.INIT_RAM_35 = 288'h30C968B45D3E57ADD6EB75BADD6CB65B2DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_36 = 288'hEB75BADD6EB75BADD6EB75BADD6EB75B6DB6AA5B64B2592C968B4510A0E4D4692D164A20;
defparam promx9_inst_14.INIT_RAM_37 = 288'hDB6D72B34AA44DE51289C4E2733CAEDBADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6;
defparam promx9_inst_14.INIT_RAM_38 = 288'hDB6DB6D96BACCD220E382C62713696DB6DD6DB75BADD6EB75BADD6EB75BADD6EB75BADB6;
defparam promx9_inst_14.INIT_RAM_39 = 288'hDB6DB2D96DB6DB6DB6CB65B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_3A = 288'hCAE56EB559A30C1ED29A556EB75CAE572D96DB65B2D96CB65B2DB6DB6DB6DB6DB65B2DB6;
defparam promx9_inst_14.INIT_RAM_3B = 288'hCB6DB2DB6CB6DB6DB6DB6572B95DB6572B95CAE56EB5489C24E134BADD72B95CAE572B95;
defparam promx9_inst_14.INIT_RAM_3C = 288'h71B8ECA0881F110A8552A954AA674940E2B279BCE6954AADD72B95CB65B2D96CB65B2D96;
defparam promx9_inst_14.INIT_RAM_3D = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6CB6572B54592194AA542A150A85429950A8533591C7E7;
defparam promx9_inst_14.INIT_RAM_3E = 288'hB31048525A2D164AA392E1F6BF6EB75BADD6CB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_14.INIT_RAM_3F = 288'hEB75BADD6EB75BADD6EB75BADD6EB75BADD6DB6DBADB6CB4D2DB0592D15C74592C968B45;

pROMX9 promx9_inst_15 (
    .DO({promx9_inst_15_dout_w[26:0],promx9_inst_15_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_31),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_15.READ_MODE = 1'b1;
defparam promx9_inst_15.BIT_WIDTH = 9;
defparam promx9_inst_15.RESET_MODE = "SYNC";
defparam promx9_inst_15.INIT_RAM_00 = 288'hDB6DB6BB5BA44DE4F2793C9E51399C4E6795DB6DBADD6EB75BADD6EB75BADD6EB75BADD6;
defparam promx9_inst_15.INIT_RAM_01 = 288'hDB6DB6DB6DB6DB6DB6CADD6A8F227A4562B168B49A4D2DAE55E554EB75BADD6DB75BADB6;
defparam promx9_inst_15.INIT_RAM_02 = 288'hDB65B6D96DB6DB2D96CAE576D95DB6DB2DB6DB6DB6DB6CB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_03 = 288'hCAE572B95CADD6EB3438B0D22F39A552EB75CAE572B95CB65B2D96CB65B2D95CAEDB2B96;
defparam promx9_inst_15.INIT_RAM_04 = 288'hCB65B6DB6CAE576D95DB6572B95CAE576DB5CAE572B95CAE56EB3474EB5E554BADD72B95;
defparam promx9_inst_15.INIT_RAM_05 = 288'h71B0F0D0361E1B8CE491A154AA552A954AA54311C6071593CE2934BAD56EB95CAE572D96;
defparam promx9_inst_15.INIT_RAM_06 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6576D96CAE56EB3422A150A8542A150A85329978923;
defparam promx9_inst_15.INIT_RAM_07 = 288'h92C99C66192D14012592D148325A2C96CFB6DB75BADD6CB65B2DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_08 = 288'hEB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADB6DB75B6DD6DB6DA698D92C168B25;
defparam promx9_inst_15.INIT_RAM_09 = 288'h99ED666F3AA551A4F279345E4F1893C9E4F2AA4CF6BB6EB6DBADD6EB75BADD6EB75BADD6;
defparam promx9_inst_15.INIT_RAM_0A = 288'hDB6DB6DB6DB6DB6DB6DB6DB2BB6CAE56EB3369038E02F48B49E4D258B49E4F26944DA4D2;
defparam promx9_inst_15.INIT_RAM_0B = 288'hDB6DB6DB6CB65B6D96CB65B2D96CAE572B95CAE572D96CB65B2BB6CB65B2DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_0C = 288'hCAE572B95CAE56EB95BADD6A93461141A534AA5D6EB75CAE572B95CB65B2D95CAE5B2DB6;
defparam promx9_inst_15.INIT_RAM_0D = 288'hCAE572D96CB65B2D96CAE572B95CAE576D95CAE572BB6CAE5B2B95CAE56E913848C2A975;
defparam promx9_inst_15.INIT_RAM_0E = 288'hF25130B2461C924AE3A2719876432A154CA552A954AA542197CE3048B4A2734AADD6EB75;
defparam promx9_inst_15.INIT_RAM_0F = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6572D96BADD6EAD132A150A8552A14C845;
defparam promx9_inst_15.INIT_RAM_10 = 288'hC6C160B258218A4A83A34968B4551C14832592C168B46DB75B6DB6CAE572DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_11 = 288'hEB75BADD6EB75B6DB6EB75BADD6EB75BADD6EB75B6DB6EB75BADD6EB75B6DD6EB6DB2B34;
defparam promx9_inst_15.INIT_RAM_12 = 288'h58B49E4F2692C5E4F279345A2F289B4562D158B4560F299E576BB6EB75BADD6EB75BADD6;
defparam promx9_inst_15.INIT_RAM_13 = 288'hCB65B2D96CB6DB2D96DB65B2DB5CB65B6B95CAED72B75AA3CD622F481C120B127A4562D1;
defparam promx9_inst_15.INIT_RAM_14 = 288'hCAE5B2DB6CAE572BB6CB65B6D96CB65B2D96CAE572B95CAE572D95CB65B2D96CAE572D96;
defparam promx9_inst_15.INIT_RAM_15 = 288'hB5C4AA975CAE572B95CADD6EB75BAD56685171ACA2734AA5D6EB95CAE572B95CB65B2B95;
defparam promx9_inst_15.INIT_RAM_16 = 288'hAA5D6EB95CAE572D96CB65B2D96DB6572B95CAE576D95CAE572B95CAE572B95CADD6A8A8;
defparam promx9_inst_15.INIT_RAM_17 = 288'h429948943B25100EE371B0DC6E392512892322A150AA552A154AA552A178B4C282C9E714;
defparam promx9_inst_15.INIT_RAM_18 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6CB6DB2D96CADD6A86742A150A85;
defparam promx9_inst_15.INIT_RAM_19 = 288'hDB6DB6D959A6364B2592C964B2582C964BC72018A4B2592C940125C3ED7ADD6CAE572DB6;
defparam promx9_inst_15.INIT_RAM_1A = 288'hEB75BADD6EB6DB6DD6EB75BADD6DB6DB6DD6DB75BADD6EB75BADD6EB75BADB6DB75B6DB6;
defparam promx9_inst_15.INIT_RAM_1B = 288'hE69C0E09037AC162D168AC5A2D27934562B058AC49EB1794CEE995DAEDB6DB6EB75BADD6;
defparam promx9_inst_15.INIT_RAM_1C = 288'hCB65B2B95CB6572B95CAE572B95CAE56EB75BA19D8D8AA9E5B2B95CADD6A9123813CE02E;
defparam promx9_inst_15.INIT_RAM_1D = 288'hCAE572B95CAE572B95CAE576D95CAE572B95CAE572BB6CAE572B95CAE5B2D95CB6572B96;
defparam promx9_inst_15.INIT_RAM_1E = 288'hCAD5266E917CD2EB75CAE572B95CADD6EB75BAD5668C238B4A6954BADD6EB75CAE572B95;
defparam promx9_inst_15.INIT_RAM_1F = 288'hE71C5A7139A556EB95CAE572B96CB6572B95CAE572B95CAE576D95CAE572B95CAE572B95;
defparam promx9_inst_15.INIT_RAM_20 = 288'h32A150A8542997896491C0DC6C361B8DC7047238E0964F22150A8542A150AA5532144D65;
defparam promx9_inst_15.INIT_RAM_21 = 288'hDAEDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB65B2D95BADD1E625;
defparam promx9_inst_15.INIT_RAM_22 = 288'hEB75BADB6DB6DB6DB6CACCF1B2592C968B24928008325A34964B05101060B0592D9F6DB6;
defparam promx9_inst_15.INIT_RAM_23 = 288'hDB6DBADD6EB75B6DD6DB75BADB6EB75BADD6DB6DB6DB6DB6DB6DB6DB6DB6DD6EB75B6DB6;
defparam promx9_inst_15.INIT_RAM_24 = 288'hAA44E67126893C5E4F071C0E090588BD629158AC49EB068BCA6774CAED76DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_25 = 288'hCAE572B95CAE572B95CADD6EB75BADD6EB75BAD52A85192B01850371205CA4EBA656EB75;
defparam promx9_inst_15.INIT_RAM_26 = 288'hCAE572B95CAE572B95CAE572B95DB6DB2B95CAE572B95CAE572B95CAE572B95CAE5B2B95;
defparam promx9_inst_15.INIT_RAM_27 = 288'hCAE572B95BAD505CEA69D52EB95CAE572B75BADD6EB75AAD5124A348BCE6954BADD6EB95;
defparam promx9_inst_15.INIT_RAM_28 = 288'h53217CB03C69416513AA556EB75CAE572B95CB6572B95CAE572B95CAE576D95CAE572B95;
defparam promx9_inst_15.INIT_RAM_29 = 288'hBAD535A4542A150A854299647A503B8D86E371B92490371B8E8965D21910A8542A150AA5;
defparam promx9_inst_15.INIT_RAM_2A = 288'h92D15E9B6CAE576DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6CB65B2B75;
defparam promx9_inst_15.INIT_RAM_2B = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB5D669AE92C164AE482C960B0582514804292C964B25;
defparam promx9_inst_15.INIT_RAM_2C = 288'hDB6DB6DB6DB6DBADD6DB75BADB6DB6DBADD6DB75BADD6EB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_2D = 288'h4141A2595CAE56EB75AA552673389B45209168B44E0906944E2733AA5D72BB5DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_2E = 288'hCAE572B95CAE572B95BADD6EB75BADD6EB75AAD56A9538A4A6C8C3B140E45028140A04C2;
defparam promx9_inst_15.INIT_RAM_2F = 288'hBADD6EB75CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B96;
defparam promx9_inst_15.INIT_RAM_30 = 288'hCAE572B95CAE572B95BAD4D91CE9A5D6EB95CAE572B95BADD6EB74AA4D187EF694D26954;
defparam promx9_inst_15.INIT_RAM_31 = 288'h42A154CA6531130903B69416514AA5D6EB75CAE572B95CAE572B95CAE572B95CAE576D95;
defparam promx9_inst_15.INIT_RAM_32 = 288'hCB65AEB75AA4D08C6543194CA853291AC92481B9186E361C91C6E3C338E47A5F2A150AA6;
defparam promx9_inst_15.INIT_RAM_33 = 288'h92C964B2592C970F95CAE576DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_34 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB2B33C6C960B2592C964B2420C17D000;
defparam promx9_inst_15.INIT_RAM_35 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DD6DB75B6DB6EB6DBADD6EB75B6DB6EB6DB6DD6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_36 = 288'h8140A05028138902C337E572B75BADD6EB74BAD52A974BA5D2E974BAE572B95CAED76DB6;
defparam promx9_inst_15.INIT_RAM_37 = 288'hCAE572B95CAE572B95CADD6EB75BADD6EB55AAD52A9349A4D2267082C11046391C8A0702;
defparam promx9_inst_15.INIT_RAM_38 = 288'h79CD2A974BADD6EB95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95;
defparam promx9_inst_15.INIT_RAM_39 = 288'hCAE572B95CAE572B95CAE572B95AAC49D270AA5D6EB95CADD6EB75BADD6EB549A4D14492;
defparam promx9_inst_15.INIT_RAM_3A = 288'h432994A85533198CA64309545C6D68C1A5349A5D6EB75CAE572B95CAE572B95CAE572B95;
defparam promx9_inst_15.INIT_RAM_3B = 288'hDB6DB2D96CADD6EB54AA4A8CD2371C08CC6532896C923B230DC6E471C0E07C671F168984;
defparam promx9_inst_15.INIT_RAM_3C = 288'h004960B2592C964B2592D168D95CAE576BB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_3D = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB59A5B60B04923948505;
defparam promx9_inst_15.INIT_RAM_3E = 288'hDB6DB2DB6DB6DB2DB6DB6DB6DB6DB6DBADD6EB75B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_15.INIT_RAM_3F = 288'h91C8A05228140A05028140A86E24030D2174BAE572D75CADD6EB95CADD72B95CAE576BB6;

pROM prom_inst_16 (
    .DO({prom_inst_16_dout_w[30:0],prom_inst_16_dout[9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_16.READ_MODE = 1'b1;
defparam prom_inst_16.BIT_WIDTH = 1;
defparam prom_inst_16.RESET_MODE = "SYNC";
defparam prom_inst_16.INIT_RAM_00 = 256'h000000000000B7FDD7FFFFFFC4000000000020C2002201208000000000000001;
defparam prom_inst_16.INIT_RAM_01 = 256'h0000CFFFFF2FFFFFE79800000500000200204000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_02 = 256'hFFC2FFFFFFE6A0400000033B9FB5FC2124000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_03 = 256'hFFFFFA001860109BEFFC579256500000000000000000000000000000000001F7;
defparam prom_inst_16.INIT_RAM_04 = 256'h13A8127E7FFFF7EB94BE00000000000000000000000000000000000FFFF203FF;
defparam prom_inst_16.INIT_RAM_05 = 256'hFDFDEFFDB2DF3A000000000000000000000000000000014FFFFE800FFFFFFFA3;
defparam prom_inst_16.INIT_RAM_06 = 256'hF265C50800000000000000000000000000000001DFFFC000BFFFFFCF380FE2EF;
defparam prom_inst_16.INIT_RAM_07 = 256'h1800000000000000000000000000000057FFF000207FFFFFFFC7B9DFFFFFDFFF;
defparam prom_inst_16.INIT_RAM_08 = 256'h0000000000000000000000000D7FE5040445FFFFEAC037BF1FFFFFFFFFDC39E0;
defparam prom_inst_16.INIT_RAM_09 = 256'h000000000000000000BFFF80510013FF3FA20396FBFFFFFFFFFEF40C9A000000;
defparam prom_inst_16.INIT_RAM_0A = 256'h000000000027FE880062004FFA7AC016FFFFFBEFFEFF6F3C6640000000000000;
defparam prom_inst_16.INIT_RAM_0B = 256'h00006FF60020000200A60C0122FFFFDFFFFFFFEAA60400000000000000000000;
defparam prom_inst_16.INIT_RAM_0C = 256'h0002040046001040401FFFF9BFFDFFFFFC6C4000010000000000000000000000;
defparam prom_inst_16.INIT_RAM_0D = 256'h110800000001FFFFDF339FDFFF7F0023000000000000000000000000000021FE;
defparam prom_inst_16.INIT_RAM_0E = 256'h00009FBFFBFEFFDFFFF06020000000800000000000000000000002AFC4004010;
defparam prom_inst_16.INIT_RAM_0F = 256'hFFFFFDEFFFFF4E004000000000000000000000000000000CE21010C842000000;
defparam prom_inst_16.INIT_RAM_10 = 256'hF77FFD90C040010000000000000000000000000320884220208800A0000007FF;
defparam prom_inst_16.INIT_RAM_11 = 256'h884000008000000000000000000000000060018400810001000000FFFFE003BF;
defparam prom_inst_16.INIT_RAM_12 = 256'h00000000000000000000000002800001000408010000003FFFF43F87FFFFFFC2;
defparam prom_inst_16.INIT_RAM_13 = 256'h00000000000000000045000410008080000000017FFF1FA43F7FCFEF40040000;
defparam prom_inst_16.INIT_RAM_14 = 256'h000000000000A00100402020088000001FFFC78DE3FFFEFFBE40800600000000;
defparam prom_inst_16.INIT_RAM_15 = 256'h0000008021410C408600000001FF79FF8917FFFFFFF014000203240000000000;
defparam prom_inst_16.INIT_RAM_16 = 256'h00400500020400000017FF1F0E00FFFFFFFF8880212440000000000000000000;
defparam prom_inst_16.INIT_RAM_17 = 256'h000880000015FFF0E10003FFFFFFF9200A009800000000000000000000001082;
defparam prom_inst_16.INIT_RAM_18 = 256'h000007EE0780000FFFFFFDE0000010C100000000000000000000000309000002;
defparam prom_inst_16.INIT_RAM_19 = 256'hE0380000BFFFFFDF000009A52100000000000000000000002002001040010000;
defparam prom_inst_16.INIT_RAM_1A = 256'h03FFE3FFF70040110240000000000000000000000020000131000480000009FF;
defparam prom_inst_16.INIT_RAM_1B = 256'hBFFB00A11040000000000000000000000000400042040808000000BFFC010000;
defparam prom_inst_16.INIT_RAM_1C = 256'h00302C000000000000000000000100000884512080000001FFF00800003FFF0B;
defparam prom_inst_16.INIT_RAM_1D = 256'h000000000000000000000804020800400950000007FF80000010FFC7DDC7D420;
defparam prom_inst_16.INIT_RAM_1E = 256'h000000000000000291C0000000090000123FC00000008FFF6FFEF03024102000;
defparam prom_inst_16.INIT_RAM_1F = 256'h000000020840800200001000000600000000003FFFFFFFD200108302A0000000;
defparam prom_inst_16.INIT_RAM_20 = 256'h48100000400101000000100000400007FEFFFFF648066741A200000000000000;
defparam prom_inst_16.INIT_RAM_21 = 256'h01500010000000000003000017FFFFFF7C804444100000000000000000000000;
defparam prom_inst_16.INIT_RAM_22 = 256'h0000000008001800007FFFFFFFC001187E889000000000000000000006340040;
defparam prom_inst_16.INIT_RAM_23 = 256'h884000400007FFFFFFA020005951082800000000000000000020409102050181;
defparam prom_inst_16.INIT_RAM_24 = 256'h00001FFFFF64E004001DC8030000000000000000000312004440410000000000;
defparam prom_inst_16.INIT_RAM_25 = 256'hFFFFF0402033CE88200000000000000000000080110002080600000000001802;
defparam prom_inst_16.INIT_RAM_26 = 256'h400031000300000000000000000000000504002000D00000000000001000087F;
defparam prom_inst_16.INIT_RAM_27 = 256'h8400000000000000000000000C400402000900000100E80040800046FFFFF380;
defparam prom_inst_16.INIT_RAM_28 = 256'h000000000020000045140100281410000000E038000400021FFFFFA4C0413F61;
defparam prom_inst_16.INIT_RAM_29 = 256'h1C08400001000810020101000004100060202000103FFFE3460013FE91428000;
defparam prom_inst_16.INIT_RAM_2A = 256'h00A40600014800100000020000C001800001FFFFEC12020209C2000000000000;
defparam prom_inst_16.INIT_RAM_2B = 256'h00008400000000400002000C000001BFFC3000013F9B80000000000000000000;
defparam prom_inst_16.INIT_RAM_2C = 256'h4000000000001000600000071DE030E10294DF60000000000000000000009801;
defparam prom_inst_16.INIT_RAM_2D = 256'h800000800300002232C40000017E6B8000000000000000000100024004282880;
defparam prom_inst_16.INIT_RAM_2E = 256'h00180000015E900000868F198000000000000000001000111019420848000010;
defparam prom_inst_16.INIT_RAM_2F = 256'h000025100C148B7AC00000000000004004200001454000150C00000000000006;
defparam prom_inst_16.INIT_RAM_30 = 256'h0840B05B0000000000000040000400010010000100000000000000002000C000;
defparam prom_inst_16.INIT_RAM_31 = 256'h72E0000000000100000000000480008010080000000000000100060006000004;
defparam prom_inst_16.INIT_RAM_32 = 256'h000000010000000000120200040100000010800000100030030000402200186E;
defparam prom_inst_16.INIT_RAM_33 = 256'h000000080000600000B0200000010800000108018000000000040044204C4000;
defparam prom_inst_16.INIT_RAM_34 = 256'h000001010500C00000001040000010800D00000000004005C28AC60000000000;
defparam prom_inst_16.INIT_RAM_35 = 256'h55440D000000008000000008005000000080000178018F800000000000000000;
defparam prom_inst_16.INIT_RAM_36 = 256'h00000008000000000007000000000000000F9C0A00000000000000000C000000;
defparam prom_inst_16.INIT_RAM_37 = 256'h410000002000200000004006408A78DB800000000000000000400000040420E0;
defparam prom_inst_16.INIT_RAM_38 = 256'h00000200000010000174C9F70000000000000000000000000089000400000000;
defparam prom_inst_16.INIT_RAM_39 = 256'h000000000002302F3C0000000000000000000000000000000000000006000000;
defparam prom_inst_16.INIT_RAM_3A = 256'h0000002283940000000000000000008000000800000000000020000000400040;
defparam prom_inst_16.INIT_RAM_3B = 256'hEEE2000000000000008000080000002104000000000104001008000600000000;
defparam prom_inst_16.INIT_RAM_3C = 256'h0000000000000000400000001480000000001800080100006000000000000A00;
defparam prom_inst_16.INIT_RAM_3D = 256'h000000000000000000500000000000820800E0000300000000000001B3E0C000;
defparam prom_inst_16.INIT_RAM_3E = 256'h00400000000000000000000000001000003800000000001185D6558000000000;
defparam prom_inst_16.INIT_RAM_3F = 256'h000000000000000060010C000001C00000000001004CC5400000000000000800;

pROM prom_inst_17 (
    .DO({prom_inst_17_dout_w[30:0],prom_inst_17_dout[9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_17.READ_MODE = 1'b1;
defparam prom_inst_17.BIT_WIDTH = 1;
defparam prom_inst_17.RESET_MODE = "SYNC";
defparam prom_inst_17.INIT_RAM_00 = 256'h0000000000C01B0000000E000001400000042E20000000000000000000080000;
defparam prom_inst_17.INIT_RAM_01 = 256'h0003F3800030007000000000000C00CE40000000000000040001800000000000;
defparam prom_inst_17.INIT_RAM_02 = 256'h000000038000000000003B9FF80000000000000020001C000000000000000000;
defparam prom_inst_17.INIT_RAM_03 = 256'h1C00000000000F4D7F4000000000000000000FE0000000000000000000000010;
defparam prom_inst_17.INIT_RAM_04 = 256'h0000401605B2C00000000000000807FC00000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_05 = 256'h677B04000000000000001FFFC000000000000000000000000000020000E00000;
defparam prom_inst_17.INIT_RAM_06 = 256'h00000000000000FE780000000000000000000000000000300003E00000000401;
defparam prom_inst_17.INIT_RAM_07 = 256'h00000000C7000000000000000000000000000000000007C800080000182BC600;
defparam prom_inst_17.INIT_RAM_08 = 256'h27E00000000000000000000000000000000000034000400210C3803C00000000;
defparam prom_inst_17.INIT_RAM_09 = 256'h0000000000000000000000000000000018000200120C93F40000000000000000;
defparam prom_inst_17.INIT_RAM_0A = 256'h00000000000000000010000000400010000080B9600000000000000001780000;
defparam prom_inst_17.INIT_RAM_0B = 256'h00000000040008000002000080380210F1000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0C = 256'h0000020000001000040100850E71000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0D = 256'h0000008000200000C1FE00000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0E = 256'h00010125050BE000000000000000000000400000000000000000000001E60020;
defparam prom_inst_17.INIT_RAM_0F = 256'h0A19FC00000000000000000000500000000000000000000001E0000000000004;
defparam prom_inst_17.INIT_RAM_10 = 256'h000000000000000000072000000000000000000007E000000000000020000801;
defparam prom_inst_17.INIT_RAM_11 = 256'h000000000000260000007FC0000000007F800000000000000100000000041420;
defparam prom_inst_17.INIT_RAM_12 = 256'h0000068000001FFF80000003F000000000000000000800000000002A00000000;
defparam prom_inst_17.INIT_RAM_13 = 256'hC00001FFFE000003C00000000000000000004000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_14 = 256'hFFF00003C00000000000000000000200000000002200000000000000000002D8;
defparam prom_inst_17.INIT_RAM_15 = 256'hC00000000000006000000010000000000280000000000000000000188C00003F;
defparam prom_inst_17.INIT_RAM_16 = 256'h30000000000000008000008004040000000000000000000035800003FFFF0001;
defparam prom_inst_17.INIT_RAM_17 = 256'hF000000004000000008000000000000000000000441000003FFFF000E0000000;
defparam prom_inst_17.INIT_RAM_18 = 256'h0020000000640A0800000000000000000602000003FFFE003000000107000000;
defparam prom_inst_17.INIT_RAM_19 = 256'h0000040000000000000000000008C000001FFFE01C0000001000000000000000;
defparam prom_inst_17.INIT_RAM_1A = 256'h0000000000000000001018000001FFFC06000000100000000000000000010000;
defparam prom_inst_17.INIT_RAM_1B = 256'h000000000000030000001FFF8180000048000000000000010000080000101401;
defparam prom_inst_17.INIT_RAM_1C = 256'h00000060000000FFE06000000400000000000000120000400000000000000000;
defparam prom_inst_17.INIT_RAM_1D = 256'h00000007FC080000090000000000000000280002000000001000000000000000;
defparam prom_inst_17.INIT_RAM_1E = 256'h7F0300000080000000000000000800001000000008800000000000000000000C;
defparam prom_inst_17.INIT_RAM_1F = 256'h0020000000000000000000000080000000040000000000000000000180000000;
defparam prom_inst_17.INIT_RAM_20 = 256'h0000000000000000000400010000000000000000000000141800000003C04000;
defparam prom_inst_17.INIT_RAM_21 = 256'h0000000000002000080008000000000000000002030000000000180000400000;
defparam prom_inst_17.INIT_RAM_22 = 256'h0000010000400210000000000000000000600000000003000014000000000000;
defparam prom_inst_17.INIT_RAM_23 = 256'h0402000000000000000000000026000000000020000100000000000000000000;
defparam prom_inst_17.INIT_RAM_24 = 256'h60000000000000000000C0000000000400014000000000000000000000000008;
defparam prom_inst_17.INIT_RAM_25 = 256'h0000000000001800000000008000000000000000000000000000000040001000;
defparam prom_inst_17.INIT_RAM_26 = 256'h0002030000000000100002000000000000000000000000000200008000000000;
defparam prom_inst_17.INIT_RAM_27 = 256'h0000000002000040000000000000000000000000001000040000000000000000;
defparam prom_inst_17.INIT_RAM_28 = 256'h0060000000000000000000000000000000008000000100000000000000000130;
defparam prom_inst_17.INIT_RAM_29 = 256'h0000000000000000000000000000040000000000000000000000000600000000;
defparam prom_inst_17.INIT_RAM_2A = 256'h000000000000000000000020000000000000000000000000C000000000040001;
defparam prom_inst_17.INIT_RAM_2B = 256'h00000000000000010000000000000000000000000C0000000000800020000000;
defparam prom_inst_17.INIT_RAM_2C = 256'h0000000008000000000000000000000209800000000010000400000000000000;
defparam prom_inst_17.INIT_RAM_2D = 256'h0040000000000000000000004030000000000300000000000000000000000000;
defparam prom_inst_17.INIT_RAM_2E = 256'h0000000000000000008700000000006000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_2F = 256'h0000000000206000000000040000000000000000000000000000000000020000;
defparam prom_inst_17.INIT_RAM_30 = 256'h00004C0000000000800020000000000000000000000000000000100000000000;
defparam prom_inst_17.INIT_RAM_31 = 256'h0000000018000800000000000000000000000000000000800000000000000000;
defparam prom_inst_17.INIT_RAM_32 = 256'h010000000000000000000000000000000000000400008000000000001FF001C0;
defparam prom_inst_17.INIT_RAM_33 = 256'h00000000000000000000000000000000200004000000000007FF801800000000;
defparam prom_inst_17.INIT_RAM_34 = 256'h000000000000000000000000010000200000000001FFF0038000000000300000;
defparam prom_inst_17.INIT_RAM_35 = 256'h00000000000000000008000000000000003FFE03700000000002000100000000;
defparam prom_inst_17.INIT_RAM_36 = 256'h0000000000004000000000000007FFC03F000000000060000000000000000000;
defparam prom_inst_17.INIT_RAM_37 = 256'h000002000000000000007FF813F8000000000400000000000000000000000000;
defparam prom_inst_17.INIT_RAM_38 = 256'h0000000000000FFC007FC000000000C000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_39 = 256'h000000FF000FFC00000000080000000000000000000000000000000000000010;
defparam prom_inst_17.INIT_RAM_3A = 256'hE200FFD000000001800000000000000000000000000000000000000080000000;
defparam prom_inst_17.INIT_RAM_3B = 256'h800000001000000000000000000070008000000000000000040000000000001F;
defparam prom_inst_17.INIT_RAM_3C = 256'h0100000000000000000003E000000000000000000020000000000001FC0007FE;
defparam prom_inst_17.INIT_RAM_3D = 256'h000000000000047FC00000000000000000010000000000003FC8007FC8000000;
defparam prom_inst_17.INIT_RAM_3E = 256'h0000009FFF00000000000000000008000000000003FC0007FC80000000300010;
defparam prom_inst_17.INIT_RAM_3F = 256'hFFFC00000000000000000040000000000063C000FFC800000002000000000000;

pROM prom_inst_18 (
    .DO({prom_inst_18_dout_w[30:0],prom_inst_18_dout[10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_18.READ_MODE = 1'b1;
defparam prom_inst_18.BIT_WIDTH = 1;
defparam prom_inst_18.RESET_MODE = "SYNC";
defparam prom_inst_18.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_18.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_02 = 256'hFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC07FF;
defparam prom_inst_18.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FFFFFFFFF;
defparam prom_inst_18.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF80383FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFC3E0F00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFF00F9C003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0B = 256'hFFFFFFFC001F8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0C = 256'h8001F80039FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0D = 256'h0E07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FE0;
defparam prom_inst_18.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDE00F0781C03FFF;
defparam prom_inst_18.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0781C01F70007FFFFFFFFF;
defparam prom_inst_18.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03E78007E0007FFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF800FE0003F000FFFFFFFFFFFFC07FFFFFFFFF;
defparam prom_inst_18.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFE0003E0007FC03DFFFFFFFFFFE003FFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_14 = 256'hFFFFFFFFFFFFC000FF801E1F071FFFFFFFFFF8121FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_15 = 256'hFFFFFF001E3E038079E1FFFFFFFFFE0070FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_16 = 256'h0780F8F001F81FFFFFFFFFE0F001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_17 = 256'h000701FFFFFFFFFF1E000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_18.INIT_RAM_18 = 256'hFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF0F003FC;
defparam prom_inst_18.INIT_RAM_19 = 256'hFFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FC000F8000F01F;
defparam prom_inst_18.INIT_RAM_1A = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0F8000CE003901FFFFFFFF;
defparam prom_inst_18.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03C003DF807103FFFFFFFFFFE0000;
defparam prom_inst_18.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE03F00703E0C107FFFFFFFFFFF00003FFFFFF;
defparam prom_inst_18.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFF033C1E00FB8108FFFFFFFFFFF80000FFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1E = 256'hFFFFFFFFFFFFFF810E3C003F01B0FFFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1F = 256'hFFFFFFFC103F0001E01E0FFFFFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_20 = 256'hB181F0003E00C0FFFFFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_21 = 256'h0E20380FFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_22 = 256'hFFFFFFFFC7FFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8C80F80;
defparam prom_inst_18.INIT_RAM_23 = 256'h0007FF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3806E01C20600;
defparam prom_inst_18.INIT_RAM_24 = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0C06383830D81FFFFFFF;
defparam prom_inst_18.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07060FE013181FFFFFF800027FC;
defparam prom_inst_18.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE06C203C01E180FFFFFF000003FE00007FF;
defparam prom_inst_18.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFF063301801C190FFFFFE0000003F00003FFFFFFFFF;
defparam prom_inst_18.INIT_RAM_28 = 256'hFFFFFFFFFFDFFFFF820B00C0100A0FFFFFC01FC003F80001FFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_29 = 256'hE3F03FFFF630700C0500C0FFFFF80FFF801FC0000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2A = 256'hFF1B01C0C0B0180FFFFF81FFFF007E00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2B = 256'h0C330381FFFFF03FFFFC07F00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1F03E3;
defparam prom_inst_18.INIT_RAM_2C = 256'h3FFFFF07FFFFE01F80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0F03C1FF8601E;
defparam prom_inst_18.INIT_RAM_2D = 256'h7FFFFF00FC0000C1FFFFFFFFFFFFFFFFFFFFFFFFFFFC0F83C0FF8181B8C61048;
defparam prom_inst_18.INIT_RAM_2E = 256'h0FE0000000FFFFFFFFFFFFFFFFFFFFFFFFE0E0FE7C0FFC0E08E6819087FFFFE0;
defparam prom_inst_18.INIT_RAM_2F = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFE0F87E3C3FFC0B883F00A01FFFFFE0FFFFFF8;
defparam prom_inst_18.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFE03C1E187FFE0CEC0E00C0FFFFFFE0FFFFFFC0FF0000;
defparam prom_inst_18.INIT_RAM_31 = 256'hFFFFFFFFFFFFFE00E00007FFF843C0600807FFFFFE0FFFFFFE07F80000000FFF;
defparam prom_inst_18.INIT_RAM_32 = 256'hFFFFFFFE0000007FFFE40C060380FFFFFFE07FFFFFE07FC00000003FFFFFFFFF;
defparam prom_inst_18.INIT_RAM_33 = 256'hF8000007FFFF807060481FFFFFFE07FFFFFE07FE00000001FFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_34 = 256'hFFFFFE06C21807FFFFFFE03FFFFFE07FF00000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_35 = 256'h223300FFFFFFFF03FFFFFE07FF800000007FFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam prom_inst_18.INIT_RAM_36 = 256'hFFFFFFF03FFFFFC0FFF800000007FFFFFFFFFFFFFFFFFFFFFFFF000003FFFFF8;
defparam prom_inst_18.INIT_RAM_37 = 256'h80FFFFF81FFFC00000003FFFFFFFFFFFFFFFFFFFFFFFF800003FFFFFE31BC01F;
defparam prom_inst_18.INIT_RAM_38 = 256'h03FFFC00000003FFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFF30780BFFFFFFFF;
defparam prom_inst_18.INIT_RAM_39 = 256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFF80000FFFFFFF0180FFFFFFFFF80FFFFF;
defparam prom_inst_18.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFF0181FFFFFFFFFC0FFFFE03FFF80;
defparam prom_inst_18.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF000007FFFFFFC083FFFFFFFFFE03FFE007FFF800000003;
defparam prom_inst_18.INIT_RAM_3C = 256'hFFFFFFFFFFF000003FFFFFFF087FFFFFFFFFE03FF000FFFF800000003FFFFFFF;
defparam prom_inst_18.INIT_RAM_3D = 256'hFFFF000003FFFFFFFC8FFFFFFFFFFF0032001FFFFC00000003FFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3E = 256'h003FFFFFFFFFFFFFFFFFFFF800000FFFFFC00000003FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFF800003FFFFFE00000003FFFFFFFFFFFFFFFFFFFFFFFFF000;

pROM prom_inst_19 (
    .DO({prom_inst_19_dout_w[30:0],prom_inst_19_dout[10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_19.READ_MODE = 1'b1;
defparam prom_inst_19.BIT_WIDTH = 1;
defparam prom_inst_19.RESET_MODE = "SYNC";
defparam prom_inst_19.INIT_RAM_00 = 256'hFFFFFFFFFF0000FFFFFFF00000003FFFFFFFFFFFFFFFFFFFFFFFFF800007FFFF;
defparam prom_inst_19.INIT_RAM_01 = 256'hFFFC007FFFFFFF80000007FFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_02 = 256'hFFFFFFFC0000007FFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_03 = 256'hE0000003FFFFFFFFFFFFFFFFFFFFFFFFFC00001FFFFFFFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_19.INIT_RAM_04 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
defparam prom_inst_19.INIT_RAM_06 = 256'hFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFF;
defparam prom_inst_19.INIT_RAM_07 = 256'hFFFFFFFC00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_08 = 256'hC01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF80000FFFFFFFFFFFFFFFFFFFFFFFFFFE07FFFF;
defparam prom_inst_19.INIT_RAM_0B = 256'hFFFFFFFFF81FFFFFFFFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0C = 256'hFE01FFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0D = 256'hFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFE01FFFF;
defparam prom_inst_19.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFE1FFFFFFFFFFFF8;
defparam prom_inst_19.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFF803FFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFC00007FF;
defparam prom_inst_19.INIT_RAM_11 = 256'hFFFFFFFFFFFF003FFFFF803FFFFFFFFF807FFFFFFFFFFFFFFE00007FFFFFFFFF;
defparam prom_inst_19.INIT_RAM_12 = 256'hFFFFF043FFFFE0007FFFFFFC0FFFFFFFFFFFFFFFFFF00003FFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_13 = 256'h3FFFFE0001FFFFFC3FFFFFFFFFFFFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_14 = 256'h000FFFFC3FFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_19.INIT_RAM_15 = 256'h3FFFFFFFFFFFFF80FFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFC103FFFFC0;
defparam prom_inst_19.INIT_RAM_16 = 256'hC00000000FFFFFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFC007FFFFC0000FFFE;
defparam prom_inst_19.INIT_RAM_17 = 256'h0FFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFF800FFFFFC0000FFF1FFFFFFF;
defparam prom_inst_19.INIT_RAM_18 = 256'hFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFF801FFFFFC0001FFCFFFFFFE00FFFFFF;
defparam prom_inst_19.INIT_RAM_19 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFF003FFFFFE0001FE3FFFFFE0FFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFE007FFFFFE0003F9FFFFFF0FFFFFFFFFFFFFFFFFFE0000;
defparam prom_inst_19.INIT_RAM_1B = 256'hFFFFFFFFFFFE00FFFFFFE0007E7FFFFF87FFFFFFFFFFFFFFFFFFF00003FFFFFF;
defparam prom_inst_19.INIT_RAM_1C = 256'hFFFFC01FFFFFFF001F9FFFFFE3FFFFFFFFFFFFFFFFFFFF80001FFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1D = 256'hFFFFFFF803F7FFFFF0FFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1E = 256'h80FCFFFFFC7FFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFF803;
defparam prom_inst_19.INIT_RAM_1F = 256'hFF1FFFFFFFFFFFFFFFFFFFFFFF00003FFFFFFFFFFFFFFFFFFFFFFF007FFFFFFF;
defparam prom_inst_19.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFF80000FFFFFFFFFFFFFFFFFFFFFFE007FFFFFFFC3FBFFF;
defparam prom_inst_19.INIT_RAM_21 = 256'hFFFFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFFE7FFFF8FFFFF;
defparam prom_inst_19.INIT_RAM_22 = 256'hFFFFFE00003FFFFFFFFFFFFFFFFFFFFFC01FFFFFFFFFFCFFFFE3FFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_23 = 256'h0001FFFFFFFFFFFFFFFFFFFFF801FFFFFFFFFFDFFFF8FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFF003FFFFFFFFFFBFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_19.INIT_RAM_25 = 256'hFFFFFFFFFFE007FFFFFFFFFF7FFFCFFFFFFFFFFFFFFFFFFFFFFFFFFF80000FFF;
defparam prom_inst_19.INIT_RAM_26 = 256'hFFFC00FFFFFFFFFFEFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFC00007FFFFFFFFF;
defparam prom_inst_19.INIT_RAM_27 = 256'hFFFFFFFFFDFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_28 = 256'hFF9FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFC00F;
defparam prom_inst_19.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000FFFFFFFFFFFFFFFFFFF801FFFFFFFF;
defparam prom_inst_19.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFC00007FFFFFFFFFFFFFFFFFF003FFFFFFFFFFBFFFC;
defparam prom_inst_19.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFE00003FFFFFFFFFFFFFFFFFE003FFFFFFFFFF7FFF9FFFFFFF;
defparam prom_inst_19.INIT_RAM_2C = 256'hFFFFFFFFF00001FFFFFFFFFFFFFFFFFC007FFFFFFFFFEFFFF3FFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2D = 256'hFF80000FFFFFFFFFFFFFFFFF800FFFFFFFFFFCFFFE7FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2E = 256'h7FFFFFFFFFFFFFFFF800FFFFFFFFFF9FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2F = 256'hFFFFFFFFFF001FFFFFFFFFFBFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000;
defparam prom_inst_19.INIT_RAM_30 = 256'hFFE003FFFFFFFFFF7FFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFF;
defparam prom_inst_19.INIT_RAM_31 = 256'hFFFFFFFFE7FFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_32 = 256'hFEFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFE00C003F;
defparam prom_inst_19.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFF8000007FFFFFFFF;
defparam prom_inst_19.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFE0000007FFFFFFFFFCFFFEF;
defparam prom_inst_19.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFC000000FFFFFFFFFFDFFFCFFFFFFFF;
defparam prom_inst_19.INIT_RAM_36 = 256'hFFFFFFFFFFFF800007FFFFFFFFF8000000FFFFFFFFFF9FFFDFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_37 = 256'hFFFFFC00003FFFFFFFFF80000007FFFFFFFFFBFFFBFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_38 = 256'h0001FFFFFFFFF00000003FFFFFFFFF3FFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_39 = 256'hFFFFFF00000001FFFFFFFFF7FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_19.INIT_RAM_3A = 256'h0000000FFFFFFFFE7FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFF;
defparam prom_inst_19.INIT_RAM_3B = 256'h7FFFFFFFEFFFEFFFFFFFFFFFFFFF8FFF7FFFFFFFFFFFFFFFF800007FFFFFFFE0;
defparam prom_inst_19.INIT_RAM_3C = 256'hFEFFFEFFFFFFFFFFFFFFF01FFFFFFFFFFFFFFFFFFFC00003FFFFFFFE00000000;
defparam prom_inst_19.INIT_RAM_3D = 256'hFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFFE00003FFFFFFFC000000007FFFFFF;
defparam prom_inst_19.INIT_RAM_3E = 256'hFFFFFF0000FFFFFFFFFFFFFFFFFFF00001FFFFFFFC000000007FFFFFFFCFFFCF;
defparam prom_inst_19.INIT_RAM_3F = 256'h0003FFFFFFFFFFFFFFFFFF80001FFFFFFF8000000007FFFFFFFDFFFDFFFFFFFF;

pROM prom_inst_20 (
    .DO({prom_inst_20_dout_w[30:0],prom_inst_20_dout[11]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_20.READ_MODE = 1'b1;
defparam prom_inst_20.BIT_WIDTH = 1;
defparam prom_inst_20.RESET_MODE = "SYNC";
defparam prom_inst_20.INIT_RAM_00 = 256'hFDFFFFFFFFF70000020000003BFFFFFFFFFFDF3DFFDDFEDF7FFFFFFFFFFFFFD2;
defparam prom_inst_20.INIT_RAM_01 = 256'hFFF20000012000001867FFFFFAFFFFFDFFDFBFFFFFFFFFFFFFFFFFFC8207EEFF;
defparam prom_inst_20.INIT_RAM_02 = 256'h0004000000195FBFFFFFFCC4604A03DEDBFFFFFFFFFFFFFFBC276FFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_03 = 256'h000005FFE79FEF641003A86DA9AFFFFFFFFFFFFFFBC0FEFFFFFFFFFFFFFFE000;
defparam prom_inst_20.INIT_RAM_04 = 256'hEC57ED81800008146B41FFFFFFFFFFFFFFFA4DFFFFFFFFFFFFFFF20000143400;
defparam prom_inst_20.INIT_RAM_05 = 256'h020210024D20C5FFFFFFFFFFFFFFF76FFFFFFFFFFFFFFA000000F3700000005C;
defparam prom_inst_20.INIT_RAM_06 = 256'h0D9A3AF7FFFFFFFFFFFFFF8FFFFFFFFFFFFFFE840000EAF8A2000030C7F01D10;
defparam prom_inst_20.INIT_RAM_07 = 256'hE7FFFFFFFFFFFFEEFFFFFFFFFFFFFFF4080005BE360000000038462000002000;
defparam prom_inst_20.INIT_RAM_08 = 256'hFFFFFFFFFBFFFFFFFFFFFFFE600000A685220000153FC800E00000000023C61F;
defparam prom_inst_20.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFE900000AA7D91A800C05DFC600000000000010BF365FFFFFF;
defparam prom_inst_20.INIT_RAM_0A = 256'hFFFFFFFFF80000A42DA242C805853FE800000410010090C399BFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0B = 256'hFF840016D893888F0359F3FEC00000200000001559FBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0C = 256'h6EE557F609FFEFBFBE000006400200000393BFFFFEFFFFFFFFFFFFFFFFFFFFFD;
defparam prom_inst_20.INIT_RAM_0D = 256'h97407FFFFFE4000020CC60200080FFDCFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_20.INIT_RAM_0E = 256'hFFFE000004010020000F9FDFFFFFFF7FFFFFFFFFFFFFFFFFFFFFB0000860D835;
defparam prom_inst_20.INIT_RAM_0F = 256'h000002100000B1FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2004B0B78927C50FFF;
defparam prom_inst_20.INIT_RAM_10 = 256'h0880026F3FBFFEFFFFFFFFFFFFFFFFFFFFFFFFE800070CCEFEEFE03FFFFFE000;
defparam prom_inst_20.INIT_RAM_11 = 256'h77BFFFFF7FFFFFFFFFFFFFFFFFFFFFEEC0A92F2FFC897F9DFFFFFE00001FEC40;
defparam prom_inst_20.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF10C14D43FFF6EE94FFFFFC0000BEC480000003D;
defparam prom_inst_20.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFF0480EB9FFE762D46FFFFFE0000D629C0803010BFFBFFFF;
defparam prom_inst_20.INIT_RAM_14 = 256'hFFFFFFFFFFF666D6BFFFC8CDF3EFFFFFC00031414C00010041BF7FF9FFFFFFFF;
defparam prom_inst_20.INIT_RAM_15 = 256'hFFFF06C56A925DFF43FEFFFFF80084AB98E80000000FEBFFFDFCDBFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_16 = 256'hA13A564FF823EFFFFF8000C19F0700000000777FDEDBBFFFFFFFFFFFFFFDFFFF;
defparam prom_inst_20.INIT_RAM_17 = 256'hFFC9FEFFFFC0000CC83E6800000006DFF5FF67FFFFFFFFFFFFFFFFFFFFFFE16C;
defparam prom_inst_20.INIT_RAM_18 = 256'hFFFE8011E4741BF00000021FFFFFEF3EFFFFFFFFFFFFFFFFFFFFFFEF688FFBDE;
defparam prom_inst_20.INIT_RAM_19 = 256'h1F272B23C0000020FFFFF65ADEFFFFFFFFFFFFFFFFFFFFBFF1BFFFF42FFF0FEF;
defparam prom_inst_20.INIT_RAM_1A = 256'h3C001C0008FFBFEEFDBFFFFFFFFFFFFFFFFFFFFF2C9E9FFE07FFDEFF7FFFE000;
defparam prom_inst_20.INIT_RAM_1B = 256'h4004FF5EEFBFFFFFFFFFFFFFFFFFFFFFFF7427FFDCFFE2C7C1FFFD0003F50154;
defparam prom_inst_20.INIT_RAM_1C = 256'hFFCBD3C20FFFFFFFFFFFFFFFFFFF43E7FF7F2EEC7007FFC0000FB8EBF9C000F4;
defparam prom_inst_20.INIT_RAM_1D = 256'h80BFFFFFFFFFFFFFFFF1E8D536A7E08B5F301FFC00007D257E7F003822382BDF;
defparam prom_inst_20.INIT_RAM_1E = 256'hFFFFFFFFFEFFFFB8B15FFF8D7DBE01FFC0003FC31434300090010FCFDBEB1FFD;
defparam prom_inst_20.INIT_RAM_1F = 256'hFFFFFFFFB0DCFFFCAFF9F00FFF4003FED16957200000002DFFEF00FD0007FFFF;
defparam prom_inst_20.INIT_RAM_20 = 256'hDAD3B7FFE4B8FEC07FF0003FF1F173DC01000009B7F9980E51881FFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_21 = 256'hFBCDDFEE03FFFFFFFFC78E11E8000000837FBB80EF19A9FFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_22 = 256'hF07FFFFD67FC6DFCDF800000003FFEC00030057FFFFFFFFFFFFFFFFFF94401FF;
defparam prom_inst_20.INIT_RAM_23 = 256'h5C33F3A2DB9C0000005FDFFC04003445FFFFFFFFFFFFFFFFFFBCC014FC6AF6FF;
defparam prom_inst_20.INIT_RAM_24 = 256'h2CA1A000009B1FF191000568DFFFFFFFFFFFFFFFFFFD3A0D7BC3AE6FCF8FFFFE;
defparam prom_inst_20.INIT_RAM_25 = 256'h00000FBF04002001DBFFFFFFFFFFFFFFFFFFF798EA197C3D7C78FFFF89CE1B97;
defparam prom_inst_20.INIT_RAM_26 = 256'hBC0080043C3FFFFFFFFFFFFFFFFFFD64E5771F8FF6938FFFD4C3CE5A8C646380;
defparam prom_inst_20.INIT_RAM_27 = 256'h1231FFFFFFFFFFFFFFFFFFF984B987FFBF7830FFB2D657FDA4E691A900000C7F;
defparam prom_inst_20.INIT_RAM_28 = 256'hFFFFFFFE3F95FFFC660D7B3FC3D73207FE35448E42279431E000005B3FA20010;
defparam prom_inst_20.INIT_RAM_29 = 256'hB1F67FFFEF5C09B7F9FF31607F84A5F99051186F9FC0001CB9FE200000B03FFF;
defparam prom_inst_20.INIT_RAM_2A = 256'hF6608EB97E67A58C0FF96240381CA8C0F05E000013EDF00472000BFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2B = 256'h0FEC79B9007F3141FE2C01041BB3FE4003CFFC140000047FFFFFFFFFFA4F27D5;
defparam prom_inst_20.INIT_RAM_2C = 256'hF81FE4A07FF88FB8E04EEDF8E21FCF008800008FFFFFFFFFFF90FB3CCFC9D002;
defparam prom_inst_20.INIT_RAM_2D = 256'hEFFFF0484748D99B6D3BFFFC200000207FFFFFFFFF18DF59D0F860607497D22F;
defparam prom_inst_20.INIT_RAM_2E = 256'h003C1B480B616FFFC00000200FFFFFFFFFF0DB7CFE4F04080DD37DCE00C1FE7C;
defparam prom_inst_20.INIT_RAM_2F = 256'hD4E5DAEFF008000018FEFFFFFFFF93B3FBC9E001780F47F2F6060E86FCFFFF81;
defparam prom_inst_20.INIT_RAM_30 = 256'hF7080200081FFFFFFFFFD0F4FCDCFC06196C13FC9E2CE0300ADFE7FC491345B4;
defparam prom_inst_20.INIT_RAM_31 = 256'h0C0B7FFFFFFFFD34E5BCF3C3BCE1811FCBE88E03882DFFFFEA1398F8E30187FB;
defparam prom_inst_20.INIT_RAM_32 = 256'hFFFFFFE9E4E9EFE073440E83F9BD01C078BD4FF7BE405CEAAD4FC23FDD808080;
defparam prom_inst_20.INIT_RAM_33 = 256'hB4EFC0100F3B00A86FA3801C0504C4FFFFE725E354A7FF9BFFFA040000039FFF;
defparam prom_inst_20.INIT_RAM_34 = 256'h81E1CA0280F2F583803C68CFFFFE76DE40D3FFFCDFFE24200C0021FFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_35 = 256'h5A59EA38380785EA7FFFE985F3C87FFFE3FFE80004000077FFFFFFFFFF5BF000;
defparam prom_inst_20.INIT_RAM_36 = 256'h0780FC3977FFFE4EDF246FFFFE27FE68104000A0B7FFFFFFFFFE7C03003E1FCA;
defparam prom_inst_20.INIT_RAM_37 = 256'hF67FFF9829F20C7FFFFB3FE0000481203DDFFFFFFFFFBF65B4A7C1FF9EB9FE7F;
defparam prom_inst_20.INIT_RAM_38 = 256'hD83F2007FFF305FE8400060003FFFFFFFFF7EF7BF61BF80FFCE883ECE0F01FE2;
defparam prom_inst_20.INIT_RAM_39 = 256'hBFFFF91FFD000000401FFFBFFFFEFFFC30240C00787600FE9C3F007E1C31FFF3;
defparam prom_inst_20.INIT_RAM_3A = 256'hFF6002900009F7FFFFFFFFFEE76A008000003E1FC007E007F9A34FFCFC37F3DF;
defparam prom_inst_20.INIT_RAM_3B = 256'h00005F7FFFFFFFF7007F3F81C00001C1F420FE01FF8A58FF39267F2FDBFFFFD5;
defparam prom_inst_20.INIT_RAM_3C = 256'hFFFFFFFD000BC1387F805C0492981FC01FFC724036B8DFFA42EFFFF06FF90000;
defparam prom_inst_20.INIT_RAM_3D = 256'hC0003BC39C783FF0332307F007FFE4CEBC4D0BFF9FBE7FFE2A7FE00000011AF7;
defparam prom_inst_20.INIT_RAM_3E = 256'h01818FFFF0C507FE00FFFF227B734D7FF929B1FB0BE7FE000020204FBFFFFFFF;
defparam prom_inst_20.INIT_RAM_3F = 256'hFFE15FFD000FFFF9D1F515DFBFDE8DD780CC7FE01C000000FBFFFFFFFA00078C;

pROM prom_inst_21 (
    .DO({prom_inst_21_dout_w[30:0],prom_inst_21_dout[11]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_21.READ_MODE = 1'b1;
defparam prom_inst_21.BIT_WIDTH = 1;
defparam prom_inst_21.RESET_MODE = "SYNC";
defparam prom_inst_21.INIT_RAM_00 = 256'hE001FFFFC98435A7F9FCB407E03467FF6000011207FFFFFFFFE0001B0037187F;
defparam prom_inst_21.INIT_RAM_01 = 256'hFF2E44E9FE0FE5888FFE367FE0003010187BFFFFFFF6001FF007598FFFFFE4BF;
defparam prom_inst_21.INIT_RAM_02 = 256'hFF003E6D28321D67FE600000008F1FFFFFFFC001C18040B1FF4C00428000BFFF;
defparam prom_inst_21.INIT_RAM_03 = 256'h7E6EC168FF800002000073FFFFFFE8003F9012CB3F000000000009FFFFF8F6FC;
defparam prom_inst_21.INIT_RAM_04 = 256'h87F98040E0010F3FFFFFFE4003C0F40533E00000000003FFFFFFF1FF1FE001F3;
defparam prom_inst_21.INIT_RAM_05 = 256'h000003FBFFFFFFFC807C23FF567E00010000003FFFFFFFE003FE200F9ACA18B7;
defparam prom_inst_21.INIT_RAM_06 = 256'h3FFFFFFDC803C71E724F80000000004FFFFFFFFFF87FE208FC4CAFC7FBFF9000;
defparam prom_inst_21.INIT_RAM_07 = 256'hFC003E73144CF80001300005FFFFFFFFFFFFFE010FE375567FEFFE200000001F;
defparam prom_inst_21.INIT_RAM_08 = 256'h2AF99C0002F3090FBFFFFFFFFFFFFFF0007F8CD93BF87FA000002043F5FFFFFF;
defparam prom_inst_21.INIT_RAM_09 = 256'h007F79FFFFFFFFFFFFFFFFFFF001FE388D05E1BFC1000800376FFFFFFED000F1;
defparam prom_inst_21.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFF5801FF071FA33DF9400000200F6FFFFFFFD400F8D1C63C0;
defparam prom_inst_21.INIT_RAM_0B = 256'hFFFFFFFFD16D01FFF065BCA63AC00400043FBFFFFFFFE4007E0FFC780007FFFE;
defparam prom_inst_21.INIT_RAM_0C = 256'hF2BEC06FFFF0A8564CE020080002F2DFFFFFFC0000FC1C3F0004FFF7FFFFFFFF;
defparam prom_inst_21.INIT_RAM_0D = 256'h9FFFE3462AFE1A381000AF1FFFF7F5C00003E80FDBE01FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0E = 256'h3E6A6000400000FBFFFF7DDCC00007FFFD7F87FFFFFFFFFFFFFFFFFFF9199E06;
defparam prom_inst_21.INIT_RAM_0F = 256'hC00000DF2FFFFFFFD8C4001FFFAD5C7FFFFFFFFFFFFFFFFECCC30FFA17FFFF9A;
defparam prom_inst_21.INIT_RAM_10 = 256'h72CFFFFFF3FE00000FFFFEC1FFFC1FFFFFFFFFFF8A4C7FFE019FFFFED376C79C;
defparam prom_inst_21.INIT_RAM_11 = 256'h8E0FB000001FCCD47FFFDEEFFFFFFDFE8E78FFFFFFFFFFFFF784A368C0304800;
defparam prom_inst_21.INIT_RAM_12 = 256'h8000EF2841FFDFF9FFFFFFF69B607FFFFFFFFED3FFF6FCE5A07400001FFBFFFB;
defparam prom_inst_21.INIT_RAM_13 = 256'h1C1FF8FFFCFFFFE433FFFFFFFFFFFFF63FFC33F92525380041FFFFFFFFFBF82F;
defparam prom_inst_21.INIT_RAM_14 = 256'hDFAFFFB733FFFFFFFFFFFF3F00FFF2B175F83008040FFBFFFFDFFFE86A001AFE;
defparam prom_inst_21.INIT_RAM_15 = 256'hFB7FFFFFFFFFF90FF387FF1CAA5B873A4000FFBFFFFFFEFD5FCA01899480FFAF;
defparam prom_inst_21.INIT_RAM_16 = 256'h2B3F3FF7CF300FFCE3D9DA0390401FF3FEFFFE7FFFBC003942781FF9FDFC7FA1;
defparam prom_inst_21.INIT_RAM_17 = 256'h89E2301FE6705FFCF4508DBF3FFFFFFFF7FE5807434D80FE9FFBE3F2347FFFF8;
defparam prom_inst_21.INIT_RAM_18 = 256'h7F7376FEFF8894877FFFFFFFFFFFFB007E7DB03FF9FEF9BC8C0FFFE0C77BE4F1;
defparam prom_inst_21.INIT_RAM_19 = 256'hB7AA2024FFFFFFFFFFFFFFE0068AB603FFAFB3C61B87FFE2C2C17A0661CF8020;
defparam prom_inst_21.INIT_RAM_1A = 256'h7FEFFFFFFFFFFFFF00C52AC07FFBF86DDFC3FF71BB0FFFEAA698A0412DFB8DF6;
defparam prom_inst_21.INIT_RAM_1B = 256'hFFFFFFFFE00D1F5807FF9FD02F88FFF8711FFFFACA6500A0082FDFB7DAEF0202;
defparam prom_inst_21.INIT_RAM_1C = 256'hF901DFFB007FFB7DC02A37F8160FFFFFC33D32744492FFFF2F5FF52087FF3FFF;
defparam prom_inst_21.INIT_RAM_1D = 256'h6007FFC7FA0F87FC16C7FFFFEA2FFCDF9B000FFC33EE7F2001BFFFFEFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1E = 256'h5EDED1BF00A0FFFFFE7BFFFF8C94103FF31DE7F80014FBBFFFFFFFFFFF503707;
defparam prom_inst_21.INIT_RAM_1F = 256'h82987FFFFF8C7FFFFF63303EFF8DC7FF8000FF7BFFFFFFFFFFF003D76C00DFED;
defparam prom_inst_21.INIT_RAM_20 = 256'hFFF11FFFFFFD1D223FE0FC7FA0000BBFBFFFDFF7FFFF807B51C04FBFBB40440F;
defparam prom_inst_21.INIT_RAM_21 = 256'hFFFFE05617FFC6067600007FF3FFFFFFFFFFF00FDF50067BFF180081F8E03FFF;
defparam prom_inst_21.INIT_RAM_22 = 256'h73DFFD4A9BD000097F3FFBBFFFFFFC01FBFB0265FFE7035074A580FFFFFE4DFF;
defparam prom_inst_21.INIT_RAM_23 = 256'hDEC780007FFBFCFEFFFFFFE01098781041F8017C134C41FFFFFFF4DFFFFFFF2D;
defparam prom_inst_21.INIT_RAM_24 = 256'h77FFB7FDEBFFFFF003D3960102FF8017C001C09AFFFFFF5BFFFFFFFF93FFFFF1;
defparam prom_inst_21.INIT_RAM_25 = 256'hFFF7EFFF00EB4EC00008564000006005F7FFFFE0FFFFFFFFF91FFFFF5CACC400;
defparam prom_inst_21.INIT_RAM_26 = 256'hFC1DB41C004180C02A00010006FFFFFC45FFFFFFFF43FFFFF86F444FE307FBFF;
defparam prom_inst_21.INIT_RAM_27 = 256'h80020058056002C0003FFFFFC17FFFFFFFFD6FFFFFC6D93BFE703F3FFFF7DAFF;
defparam prom_inst_21.INIT_RAM_28 = 256'h00F000540004FF7FF807FFFFFFFFA53FFFFE204137FF8573EE7E7FFFFC019FF5;
defparam prom_inst_21.INIT_RAM_29 = 256'h00000FFFFF061FFFFFFFFF0FFFFFF1F7B0FFF953FFEFF75EFE40377BB8000000;
defparam prom_inst_21.INIT_RAM_2A = 256'hFF7E0DFFFFFFFFD55FFFFF8DACDDFFE73F6A39E3F782069383000000000A800F;
defparam prom_inst_21.INIT_RAM_2B = 256'hFFFFFFFE1BFFFFFD6ABCBBFDF3E774F7D39000CE1D700000000270016800011F;
defparam prom_inst_21.INIT_RAM_2C = 256'hF83FFFFFE3295CFFE75E7FEE033A003B1EEE000000006E00270000017DFFE44F;
defparam prom_inst_21.INIT_RAM_2D = 256'hFF304A43FC13FBDB1C00001F5C68E0000000040007B0000086FFF839FFFFFFFF;
defparam prom_inst_21.INIT_RAM_2E = 256'h1FFF3FF7EF1E8003CE645C00000000B400FA000004A3FFC2AFFFFFFFFF2BFFFF;
defparam prom_inst_21.INIT_RAM_2F = 256'hFF910001E0FBF9C000000018800BE0000000DFFF28FFFFFFFFF51FFFFFF9B0C0;
defparam prom_inst_21.INIT_RAM_30 = 256'h38D3363C000000013001CC0000004CE5F403FFFFFFFF5FFFFFFF941243FDF3FC;
defparam prom_inst_21.INIT_RAM_31 = 256'h8000000037002CC000000000FF8EDFFFFFFFF5DFFFFFFC6A2A77CFFFE6DE4004;
defparam prom_inst_21.INIT_RAM_32 = 256'h04200778000000000FEC417FFFFFFE87FFFFFFE750405FF0FFDDC00034E0D813;
defparam prom_inst_21.INIT_RAM_33 = 256'h8000000003FEB3C3FFFFFFE1FFFFFFFFF8700AFFAFFE6200040D399D38000000;
defparam prom_inst_21.INIT_RAM_34 = 256'h0801FE0EBFFFFFFDFFFFFFFFFDA42C7FF364BFA40381F57E31800000006600D9;
defparam prom_inst_21.INIT_RAM_35 = 256'hB97FFFFF37FFFFFFFFEC0089FF1D7FC000501FDDEB3C00000009400D38000000;
defparam prom_inst_21.INIT_RAM_36 = 256'h9DB7FFFFFFFEE3128FF10FE4000C03A89691C0000001D801CF000000000009B8;
defparam prom_inst_21.INIT_RAM_37 = 256'hFFFFF340F04F71D0810101F91F1CDC0000001D803560000000000017874FFFFF;
defparam prom_inst_21.INIT_RAM_38 = 256'h7267F0003C00083ACEE084C0000002B0034E0000000000001067D9FF300EFFFF;
defparam prom_inst_21.INIT_RAM_39 = 256'h3F500F83AA9E014E0000002F00EEE00000000000000158EAEC085FFFFFFFFF48;
defparam prom_inst_21.INIT_RAM_3A = 256'h6EFD607AE0000004B00D8C000000000000000996840AA9FFFFFFFFF843714F00;
defparam prom_inst_21.INIT_RAM_3B = 256'hA6000000BA01D5E0000000000006186157E7D47FFFFFFFFFCD8481F001C00060;
defparam prom_inst_21.INIT_RAM_3C = 256'h04E01D1E00000000004FE0A1A0FFD20FFFFFFFFEEA6189450086000F8F3E1E02;
defparam prom_inst_21.INIT_RAM_3D = 256'hC0000000001FEC7EC1F7178FFFFFFFFFFECE1210400040003D878DE00EF00000;
defparam prom_inst_21.INIT_RAM_3E = 256'h000FF18FFDC3E003FFFFFFFFFFFC4802830002001CFE5B4C254E0000001401AB;
defparam prom_inst_21.INIT_RAM_3F = 256'hFFF5A401DDFFFFFFFFFFFE84C000000007A1849406367000000AC018BE000000;

pROM prom_inst_22 (
    .DO({prom_inst_22_dout_w[30:0],prom_inst_22_dout[12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_22.READ_MODE = 1'b1;
defparam prom_inst_22.BIT_WIDTH = 1;
defparam prom_inst_22.RESET_MODE = "SYNC";
defparam prom_inst_22.INIT_RAM_00 = 256'hFFFFFFFFFFF70000020000003BFFFFFFFFFFDF3DFFDDFEDF7FFFFFFFFFFFFFFD;
defparam prom_inst_22.INIT_RAM_01 = 256'hFFF20000012000001867FFFFFAFFFFFDFFDFBFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_02 = 256'h001C000000195FBFFFFFFCC4604A03DEDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_03 = 256'h000005FFE79FEF641003A86DA9AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_22.INIT_RAM_04 = 256'hEC57ED81800008146B41FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2000014F000;
defparam prom_inst_22.INIT_RAM_05 = 256'h020210024D20C5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0000007FD00000005C;
defparam prom_inst_22.INIT_RAM_06 = 256'h0D9A3AF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE840000FFFFE2000030C7F01D10;
defparam prom_inst_22.INIT_RAM_07 = 256'hE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF4080004FFDB0000000038462000002000;
defparam prom_inst_22.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE600001E3F9BE0000153FC800E00000000023C61F;
defparam prom_inst_22.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFE9000009F4EBFF800C05DFC600000000000010BF365FFFFFF;
defparam prom_inst_22.INIT_RAM_0A = 256'hFFFFFFFFF80000A7F92DFF8805853FE800000410010090C399BFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0B = 256'hFF840017FFE2FFFF0359F3FEC00000200000001559FBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0C = 256'h3FFF73FFDBFFEFBFBE000006400200000393BFFFFEFFFFFFFFFFFFFFFFFFFFFD;
defparam prom_inst_22.INIT_RAM_0D = 256'hE0F87FFFFFE4000020CC60200080FFDCFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_22.INIT_RAM_0E = 256'hFFFE000004010020000F9FDFFFFFFF7FFFFFFFFFFFFFFFFFFFFFB0001BFF938F;
defparam prom_inst_22.INIT_RAM_0F = 256'h000002100000B1FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2007EFE77FBFBFEFFF;
defparam prom_inst_22.INIT_RAM_10 = 256'h0880026F3FBFFEFFFFFFFFFFFFFFFFFFFFFFFFE8007B7EBFAC37FFBFFFFFE000;
defparam prom_inst_22.INIT_RAM_11 = 256'h77BFFFFF7FFFFFFFFFFFFFFFFFFFFFEEC0BFEE3BFF6EFFF7FFFFFE00001F9C40;
defparam prom_inst_22.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF103FFBF7FFA07FE5FFFFFC0000BB3480000003D;
defparam prom_inst_22.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFF04FFFE0FFFEEBF9AFFFFFE0000C99FC0803010BFFBFFFF;
defparam prom_inst_22.INIT_RAM_14 = 256'hFFFFFFFFFFF65FFFAF3FEDE5FAEFFFFFC0003ED59C00010041BF7FF9FFFFFFFF;
defparam prom_inst_22.INIT_RAM_15 = 256'hFFFF027FCFC9FD7F75FEFFFFF800874890E80000000FEBFFFDFCDBFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_16 = 256'h7BFF1B67FE6BEFFFFF8000ED667500000000777FDEDBBFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_17 = 256'hFFECFEFFFFC0000FF05FE800000006DFF5FF67FFFFFFFFFFFFFFFFFFFFFFE11C;
defparam prom_inst_22.INIT_RAM_18 = 256'hFFFE8011FF8FFF700000021FFFFFEF3EFFFFFFFFFFFFFFFFFFFFFFECA7A7FCDA;
defparam prom_inst_22.INIT_RAM_19 = 256'h1FF3FFBFC0000020FFFFF65ADEFFFFFFFFFFFFFFFFFFFFBFE6BBFFF3BFFE5FEF;
defparam prom_inst_22.INIT_RAM_1A = 256'h7C001C0008FFBFEEFDBFFFFFFFFFFFFFFFFFFFFF2C03FFFFCCFFD77EFFFFE000;
defparam prom_inst_22.INIT_RAM_1B = 256'h4004FF5EEFBFFFFFFFFFFFFFFFFFFFFFFF6027FFD593F8FFDFFFFD0003FBFFDC;
defparam prom_inst_22.INIT_RAM_1C = 256'hFFCBD3C20FFFFFFFFFFFFFFFFFFF076FF6F88FBD7DFFFFC0000FD7E765C000F4;
defparam prom_inst_22.INIT_RAM_1D = 256'h80BFFFFFFFFFFFFFFFF1F02D7EDFF71FC6AFFFFC00007EF9645F003822382BDF;
defparam prom_inst_22.INIT_RAM_1E = 256'hFFFFFFFFFEFFFFC38D97FFD6FC16FFFFC0003FF1CA0A300090010FCFDBEB1FFD;
defparam prom_inst_22.INIT_RAM_1F = 256'hFFFFFFFE187F7FFEEFEFFFFFFF4003FF4A96AB200000002DFFEF00FD0007FFFF;
defparam prom_inst_22.INIT_RAM_20 = 256'hD40077FFBBFDBF3FFFF0003FFD0E421C01000009B7F9980E51881FFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_21 = 256'hFDFFCFE1FFFFFFFFFFF7712EE8000000837FBB80EF19A9FFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_22 = 256'h0FFFFFFA87FFAD31E7800000003FFEC00030057FFFFFFFFFFFFFFFFFF8DC0BFF;
defparam prom_inst_22.INIT_RAM_23 = 256'hDD1BFD2D847C0000005FDFFC04003445FFFFFFFFFFFFFFFFFFC2C085FED9FAFE;
defparam prom_inst_22.INIT_RAM_24 = 256'h539EA000009B1FF191000568DFFFFFFFFFFFFFFFFFFE1C065FB78EA7E07FFFFF;
defparam prom_inst_22.INIT_RAM_25 = 256'h00000FBF04002001DBFFFFFFFFFFFFFFFFFFE0407855F914F807FFFF5D0B5FE1;
defparam prom_inst_22.INIT_RAM_26 = 256'hBC0080043C3FFFFFFFFFFFFFFFFFFE098071BF9AEEC07FFFE63FBA7F2F9F9380;
defparam prom_inst_22.INIT_RAM_27 = 256'h1231FFFFFFFFFFFFFFFFFFE0146987FFBEC10FFFBFBF5F93B979AE2900000C7F;
defparam prom_inst_22.INIT_RAM_28 = 256'hFFFFFFFFFFB5FFFF41157A7FC7D921FFFFF7AF17BBCBC3CFE000005B3FA20010;
defparam prom_inst_22.INIT_RAM_29 = 256'hEDF2BFFFFE2CF1B7FDFE701FFFF26401433E7F91BFC0001CB9FE200000B03FFF;
defparam prom_inst_22.INIT_RAM_2A = 256'hFFB902587FD79D93FFFE7B3FC2D4F3F72F7E000013EDF00472000BFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2B = 256'h0F9D7A7BFFFFDB2FFFC94FDFFC2BFE4003CFFC140000047FFFFFFFFFFE6FBBD9;
defparam prom_inst_22.INIT_RAM_2C = 256'hA7FFF8BDFFFF342EFDF85FF8E21FCF008800008FFFFFFFFFFFDFFCFEFFF0E800;
defparam prom_inst_22.INIT_RAM_2D = 256'hDFFFFD3DF7B742D4ED3BFFFC200000207FFFFFFFFF1F2F41FFFF82408431E2F3;
defparam prom_inst_22.INIT_RAM_2E = 256'hDFBBF04003E16FFFC00000200FFFFFFFFFE2E47D7D3FF8120893FC5F083FFFBE;
defparam prom_inst_22.INIT_RAM_2F = 256'hEFE7DAEFF008000018FFFFFFFFFFE7C7E7F1FFE1ED0A77D8E001FFFBA3FFFFEF;
defparam prom_inst_22.INIT_RAM_30 = 256'hF7080200081FFFFFFFFFFF7D3D397FF900B407FD7E0C1FFFBEBFE7FF7F7D7810;
defparam prom_inst_22.INIT_RAM_31 = 256'h0C0B7FFFFFFFFFC0F8600FFC3C8041BFFFE881FFF0EBFFFFF0DFE90275FF87FB;
defparam prom_inst_22.INIT_RAM_32 = 256'hFFFFFFFD0106007F83EA1283FB3C003FFF15BFF7BFBFBF614E7FFE7FDD808080;
defparam prom_inst_22.INIT_RAM_33 = 256'hB3100007F03FA0307FD38003FFFA53FFFFFA7BFB06FFFFF9FFFA040000039FFF;
defparam prom_inst_22.INIT_RAM_34 = 256'h7E01FA0200CBF9807FFFBFFFFFFFACBF9DDFFFFFCFFE24200C0021FFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_35 = 256'h174EEEB807FFF88DFFFFF353FD09FFFFFCFFE80004000077FFFFFFFFFFE40000;
defparam prom_inst_22.INIT_RAM_36 = 256'h007FFFDAAFFFFF3EBFCCFFFFFFE3FE68104000A0BFFFFFFFFFFF800383C01FC6;
defparam prom_inst_22.INIT_RAM_37 = 256'h6EFFFFEA47FCAFFFFFFF3FE0000481203DFFFFFFFFFFF875C79801FF8A895E5F;
defparam prom_inst_22.INIT_RAM_38 = 256'hECFFC8FFFFFFE7FE8400060003FFFFFFFFFFFFFCC6E4000FFCB043E4E00FFFFC;
defparam prom_inst_22.INIT_RAM_39 = 256'hFFFFFF1FFD000000401FFFFFFFFFFFFFB01FF0007871027F1C00FFFFEED7FFFD;
defparam prom_inst_22.INIT_RAM_3A = 256'hFF6002900009FFFFFFFFFFFFF7EBFE800000021FD0001FFFFE6EBFFF792FFD5F;
defparam prom_inst_22.INIT_RAM_3B = 256'h00005FFFFFFFFFFFFF7FFFF1C0000061F42001FFFFF03FFFCEFDFFC6FFFFFFF7;
defparam prom_inst_22.INIT_RAM_3C = 256'hFFFFFFFFFFFFC43FFF8000050298003FFFFFBF5FCFA4BFFCC7FFFFFF7FF90000;
defparam prom_inst_22.INIT_RAM_3D = 256'hFFFFF863F7F800003043000FFFFFF9F3C7F377FFE8FFFFFFE1FFE00000011AFF;
defparam prom_inst_22.INIT_RAM_3E = 256'hFF7F800000C60001FFFFFFC3D0EED4FFFE67FFFFFEDFFE000020204FFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3F = 256'h0000E002FFFFFFFEFFCFE13FBFE5BFFFFFCFFFE01C000000FFFFFFFFFFFFFF86;

pROM prom_inst_23 (
    .DO({prom_inst_23_dout_w[30:0],prom_inst_23_dout[12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_23.READ_MODE = 1'b1;
defparam prom_inst_23.BIT_WIDTH = 1;
defparam prom_inst_23.RESET_MODE = "SYNC";
defparam prom_inst_23.INIT_RAM_00 = 256'h1FFFFFFFF29FEB9FF9FF2DFFFFF01FFF6000011207FFFFFFFFFFFF79FFF0F800;
defparam prom_inst_23.INIT_RAM_01 = 256'hFFC85DA7FE0FF96FFFFE01FFE0003010187FFFFFFFFFFFE59FFE078000001F40;
defparam prom_inst_23.INIT_RAM_02 = 256'hFF003F8B7FF3FD9FFE600000008FFFFFFFFFFFFE41FFF07000B3FFFD7FFFFFFF;
defparam prom_inst_23.INIT_RAM_03 = 256'h5BFEFF67FF80000200007FFFFFFFFFFFC31FF3C700FFFFFFFFFFFFFFFFFF3F1B;
defparam prom_inst_23.INIT_RAM_04 = 256'h5FF98040E0010FFFFFFFFFFFFC04F41CF01FFFFFFFFFFFFFFFFFFE00FFE001FC;
defparam prom_inst_23.INIT_RAM_05 = 256'h000003FFFFFFFFFFFF802806CE01FFFFFFFFFFFFFFFFFFFFFFFE200FE3BF1F40;
defparam prom_inst_23.INIT_RAM_06 = 256'hFFFFFFFFFFFC07A1C9C07FFFFFFFFFFFFFFFFFFFFFFFE208FF8ADFFC05FF9000;
defparam prom_inst_23.INIT_RAM_07 = 256'hFFFFC07ED93C07FFFFFFFFFFFFFFFFFFFFFFFE010FFC667D8057FE200000001F;
defparam prom_inst_23.INIT_RAM_08 = 256'hC76783FFFFFFFFFFFFFFFFFFFFFFFFF0007FF0E27403BFA000002043FFFFFFFF;
defparam prom_inst_23.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF001FFC0EEE307BFC100080037FFFFFFFFFFFF01;
defparam prom_inst_23.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFF801FFF81374F3F9400000200FFFFFFFFFFFFF00C7BE03F;
defparam prom_inst_23.INIT_RAM_0B = 256'hFFFFFFFFE7FD01FFFF87C2D3BAC00400043FFFFFFFFFFFFF800FFC07FFFFFFFF;
defparam prom_inst_23.INIT_RAM_0C = 256'hFFFDC06FFFFF3BA8BCE020080002FFFFFFFFFFFFFF001C00FFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0D = 256'h9FFFFDD905BE1A381000AFFFFFFFFFFFFFFC0000241FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0E = 256'hE9146000400000FFFFFFFFFFFFFFF80000807FFFFFFFFFFFFFFFFFFFFDBB7E06;
defparam prom_inst_23.INIT_RAM_0F = 256'hC00000DFFFFFFFFFFFFFFFE0007703FFFFFFFFFFFFFFFFFFFAF8FFFA17FFFFEE;
defparam prom_inst_23.INIT_RAM_10 = 256'h7FFFFFFFFFFFFFFFF000FA3FFFFFFFFFFFFFFFFFEFCBFFFE019FFFFF74A1179C;
defparam prom_inst_23.INIT_RAM_11 = 256'hFFFFFFFFFFE1DEB3FFFF9E5FFFFFFDFDDE57FFFFFFFFFFFFFB3014A8C0304800;
defparam prom_inst_23.INIT_RAM_12 = 256'hFFFF1F993FFFFFFFBFFFFFFBBF1FFFFFFFFFFED3FFD90013A07400001FFFFFFF;
defparam prom_inst_23.INIT_RAM_13 = 256'h53FFFDFFFDFFFFFE2FFFFFFFFFFFFFF63FFF4E44D525380041FFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_14 = 256'hFFEFFFFF2FFFFFFFFFFFFFFF00FFFB4E8A783008040FFFFFFFFFFFFFFFFFE1EF;
defparam prom_inst_23.INIT_RAM_15 = 256'h97FFFFFFFFFFFEE77387FFDB11C7873A4000FFFFFFFFFFFFFFFFFE38F67FFFFF;
defparam prom_inst_23.INIT_RAM_16 = 256'hAFFFFFFFC7300FFEDC12BA0390401FFFFFFFFFFFFFFFFFC01BA7FFFDFFFFFFFF;
defparam prom_inst_23.INIT_RAM_17 = 256'h24E2301FF78D11FCF4508DBFFFFFFFFFFFFFFFF841747FFFDFFFEFFE7BFFFFFF;
defparam prom_inst_23.INIT_RAM_18 = 256'h7FBE010EFF889487FFFFFFFFFFFFFFFF8B3A8FFFFDFFFDFF39FFFFFCF13BFB1E;
defparam prom_inst_23.INIT_RAM_19 = 256'h77AA2024FFFFFFFFFFFFFFFFF802D1FFFFFFFFFFE97FFFFCD63FFFE667BF8020;
defparam prom_inst_23.INIT_RAM_1A = 256'h7FFFFFFFFFFFFFFFFF104E3FFFFDFFFBF77FFFFED0FFFFEA260038412DFDF3CC;
defparam prom_inst_23.INIT_RAM_1B = 256'hFFFFFFFFFFF17DC7FFFFFFFE79A7FFFFFCFFFFFE02250020082FEEB807EF0202;
defparam prom_inst_23.INIT_RAM_1C = 256'hFFFE5DA8FFFFFE7FDFE1FFFFC8FFFFFF830136480492FF70383FF52087FFFFFF;
defparam prom_inst_23.INIT_RAM_1D = 256'h1FFFFFFFFDED7FFFEFBFFFFFF01FFFE403000FF8F011FF2001BFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1E = 256'hBEFB4FFFFD5FFFFFFF07FFFFEC14103FD42C07F80014FFFFFFFFFFFFFFFFC135;
defparam prom_inst_23.INIT_RAM_1F = 256'hFDF7FFFFFFE0FFFFFFA0303EFEB0461F8000FFFFFFFFFFFFFFFFFC46A3FFFFFF;
defparam prom_inst_23.INIT_RAM_20 = 256'hFFFC8FFFFFFE01223FF94000A0000BBFFFFFFFFFFFFFFF83C43FFFFFFD7F73FF;
defparam prom_inst_23.INIT_RAM_21 = 256'hFFFFF02E17FF88C08600007FFFFFFFFFFFFFFFF3E5CFFFFFFFE7E67FFF73FFFF;
defparam prom_inst_23.INIT_RAM_22 = 256'hF3DFFF10285000097FFFFFFFFFFFFFFE6FE8FFFFFFFFFDCFFFCA7FFFFFFF83FF;
defparam prom_inst_23.INIT_RAM_23 = 256'h0F0180007FFFFFFFFFFFFFFFE0FD07FFFFFFFFABFFF63FFFFFFFF83FFFFFFFD0;
defparam prom_inst_23.INIT_RAM_24 = 256'h77FFFFFFFFFFFFFFFCD731FFFFFFFFE93FFFDFFFFFFFFF83FFFFFFFE87FFFFE2;
defparam prom_inst_23.INIT_RAM_25 = 256'hFFFFFFFFFF0BAA3FFFFFFFFE8FFFA7FFFFFFFFF83FFFFFFFF09FFFFF80822400;
defparam prom_inst_23.INIT_RAM_26 = 256'hFFE33743FFFFFFFFD5FFF6FFFFFFFFFF83FFFFFFFFC3FFFFFC85804FE307FFFF;
defparam prom_inst_23.INIT_RAM_27 = 256'h7FFFFFFFFA9FFDFFFFFFFFFFF83FFFFFFFFB0FFFFFE180C3FE703FFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_28 = 256'hFF27FFB3FFFFFFFFFF03FFFFFFFFC2BFFFFF001037FF85FFFFFFFFFFFFFE7D9C;
defparam prom_inst_23.INIT_RAM_29 = 256'h7FFFFFFFFFF63FFFFFFFFD0FFFFFF80613FFF95FFFFFFFFFFFFFC6BA87FFFFFF;
defparam prom_inst_23.INIT_RAM_2A = 256'hFFFF81FFFFFFFFEC1FFFFFC0881DFFE7FFFFFFFFFFFFF891D0FFFFFFFFF07FF7;
defparam prom_inst_23.INIT_RAM_2B = 256'hFFFFFFFF03FFFFFF03C03BFDFFFFFFFFFFFFFF0F370FFFFFFFFD2FFE67FFFFFF;
defparam prom_inst_23.INIT_RAM_2C = 256'hF03FFFFFF00060FFE7FFFFFFFFFFFFC126A1FFFFFFFF9DFFCAFFFFFFFFFFF81F;
defparam prom_inst_23.INIT_RAM_2D = 256'hFFE05047FC1FFFFFFFFFFFE05A741FFFFFFFFABFF94FFFFFFFFFFFF8FFFFFFFF;
defparam prom_inst_23.INIT_RAM_2E = 256'h1FFFFFFFFFFFFFFC060AC3FFFFFFFF43FF11FFFFFFFFFFFC87FFFFFFFFA3FFFF;
defparam prom_inst_23.INIT_RAM_2F = 256'hFFFFFFFE01D9283FFFFFFFE87FF29FFFFFFFFFFFC87FFFFFFFF8DFFFFFFD3418;
defparam prom_inst_23.INIT_RAM_30 = 256'hC0EBF503FFFFFFFEEFFE33FFFFFFFFFFFE03FFFFFFFF81FFFFFFE00703FDFFFF;
defparam prom_inst_23.INIT_RAM_31 = 256'h7FFFFFFFD8FFC23FFFFFFFFFFFF61FFFFFFFF83FFFFFFF40200FCFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_32 = 256'hF91FF9A7FFFFFFFFFFFF80FFFFFFFF1BFFFFFFFA01427FFFFFFFFFFFF33FFFB0;
defparam prom_inst_23.INIT_RAM_33 = 256'h7FFFFFFFFFFFFFC3FFFFFFF43FFFFFFF905C83FFFFFFFFFFFFF2346B07FFFFFF;
defparam prom_inst_23.INIT_RAM_34 = 256'hFFFFFFEE3FFFFFFE07FFFFFFFE843C3FFFFFFFFFFC7E056F707FFFFFFFB9FF14;
defparam prom_inst_23.INIT_RAM_35 = 256'h79FFFFFFC07FFFFFFFF40187FFFFFFFFFF8FE2FFD703FFFFFFF43FF287FFFFFF;
defparam prom_inst_23.INIT_RAM_36 = 256'hE00FFFFFFFFF23510FFFFFFFFFF3FC28AA703FFFFFFE57FE78FFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_37 = 256'hFFFFFD20C06FFFFFFFFE7E0924EBC3FFFFFFE47FC51FFFFFFFFFFFFFFACFFFFF;
defparam prom_inst_23.INIT_RAM_38 = 256'h3043FFFFFFFFEFC26E9F1C3FFFFFFCAFFCE1FFFFFFFFFFFFFF8FDCFFF801FFFF;
defparam prom_inst_23.INIT_RAM_39 = 256'hFFFFF07C1819FAC1FFFFFFD8FF0A1FFFFFFFFFFFFFFE28EA4000BFFFFFFFFFE8;
defparam prom_inst_23.INIT_RAM_3A = 256'hB2F31FA61FFFFFF84FF0C3FFFFFFFFFFFFFFF0FE8402A7FFFFFFFFFF4F511FFF;
defparam prom_inst_23.INIT_RAM_3B = 256'hE1FFFFFF79FE1C1FFFFFFFFFFFF9CF8E7FE7F3FFFFFFFFFFF20542FFFFFFFF9F;
defparam prom_inst_23.INIT_RAM_3C = 256'hF99FE381FFFFFFFFFFB01BCE077BF1FFFFFFFFFFFF9108C7FFFFFFF1707E21FD;
defparam prom_inst_23.INIT_RAM_3D = 256'h3FFFFFFFFFE005FF3E07307FFFFFFFFFFFFD82001FFFFFFF821F889FCA0FFFFF;
defparam prom_inst_23.INIT_RAM_3E = 256'hFFF0016FFE3C1FFFFFFFFFFFFFFFF41283FFFFFFE284DB93F8A1FFFFFFA3FE28;
defparam prom_inst_23.INIT_RAM_3F = 256'hFFF85BFFFFFFFFFFFFFFFF26C01FFFFFF82444917FFA0FFFFFF63FE381FFFFFF;

pROM prom_inst_24 (
    .DO({prom_inst_24_dout_w[30:0],prom_inst_24_dout[13]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_24.READ_MODE = 1'b1;
defparam prom_inst_24.BIT_WIDTH = 1;
defparam prom_inst_24.RESET_MODE = "SYNC";
defparam prom_inst_24.INIT_RAM_00 = 256'hFFFFFFFFFFF70000020000003BFFFFFFFFFFDF3DFFDDFEDF7FFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_01 = 256'hFFF20000012000001867FFFFFAFFFFFDFFDFBFFFFFFFFFFFFFFFFFFFEFFFFFFF;
defparam prom_inst_24.INIT_RAM_02 = 256'h001E000000195FBFFFFFFCC4604A03DEDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_03 = 256'h000005FFE79FEF641003A86DA9AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_24.INIT_RAM_04 = 256'hEC57ED81800008146B41FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2000016F800;
defparam prom_inst_24.INIT_RAM_05 = 256'h020210024D20C5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA000000FFF00000005C;
defparam prom_inst_24.INIT_RAM_06 = 256'h0D9A3AF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE840000FFFF62000030C7F01D10;
defparam prom_inst_24.INIT_RAM_07 = 256'hE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF4080005FFFF0000000038462000002000;
defparam prom_inst_24.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE600001E7FDFE0000153FC800E00000000023C61F;
defparam prom_inst_24.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFE900000BF5FBFF800C05DFC600000000000010BF365FFFFFF;
defparam prom_inst_24.INIT_RAM_0A = 256'hFFFFFFFFF80000AFFD6FFFC805853FE800000410010090C399BFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0B = 256'hFF840017FFF3FFFD0359F3FEC00000200000001559FBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0C = 256'h7FFF17FFDFFFEFBFBE000006400200000393BFFFFEFFFFFFFFFFFFFFFFFFFFFD;
defparam prom_inst_24.INIT_RAM_0D = 256'hF3F87FFFFFE4000020CC60200080FFDCFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_24.INIT_RAM_0E = 256'hFFFE000004010020000F9FDFFFFFFF7FFFFFFFFFFFFFFFFFFFFFB0001FFFDB9F;
defparam prom_inst_24.INIT_RAM_0F = 256'h000002100000B1FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2007FFF7FF7FFFEFFF;
defparam prom_inst_24.INIT_RAM_10 = 256'h0880026F3FBFFEFFFFFFFFFFFFFFFFFFFFFFFFE800FF7EFFFCBFFFBFFFFFE000;
defparam prom_inst_24.INIT_RAM_11 = 256'h77BFFFFF7FFFFFFFFFFFFFFFFFFFFFEEC0BFFFBFFFEFFFFFFFFFFE00001FFC40;
defparam prom_inst_24.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF107FFFF7FFFCFFF7FFFFFC0000BE0C80000003D;
defparam prom_inst_24.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFF05FFFBDFFFFEBFD9FFFFFE0000F11BC0803010BFFBFFFF;
defparam prom_inst_24.INIT_RAM_14 = 256'hFFFFFFFFFFF67FFFBB7FEDEDFB1FFFFFC000304D3C00010041BF7FF9FFFFFFFF;
defparam prom_inst_24.INIT_RAM_15 = 256'hFFFF06FFEFD9FDFFF7C1FFFFF8008707E0E80000000FEBFFFDFCDBFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_16 = 256'hFBFF576FFEEC1FFFFF8000F30E5B00000000777FDEDBBFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_17 = 256'hFFE701FFFFC0000E0E501800000006DFF5FF67FFFFFFFFFFFFFFFFFFFFFFE11E;
defparam prom_inst_24.INIT_RAM_18 = 256'hFFFE8011F08000F00000021FFFFFEF3EFFFFFFFFFFFFFFFFFFFFFFEF6FAFFDDE;
defparam prom_inst_24.INIT_RAM_19 = 256'h1F88006FC0000020FFFFF65ADEFFFFFFFFFFFFFFFFFFFFBFFDBFFFF7FFFF681F;
defparam prom_inst_24.INIT_RAM_1A = 256'h7C001C0008FFBFEEFDBFFFFFFFFFFFFFFFFFFFFF2FF7FFFFCDFFDA01FFFFE000;
defparam prom_inst_24.INIT_RAM_1B = 256'h4004FF5EEFBFFFFFFFFFFFFFFFFFFFFFFF7FD7FFDEF7FB201FFFFD0003FC002C;
defparam prom_inst_24.INIT_RAM_1C = 256'hFFCBD3C20FFFFFFFFFFFFFFFFFFEFCEFFFFD9FE28AFFFFC0000FEC17E3C000F4;
defparam prom_inst_24.INIT_RAM_1D = 256'h80BFFFFFFFFFFFFFFFF1FFCB7EFFF754291FFFFC00007F47254F003822382BDF;
defparam prom_inst_24.INIT_RAM_1E = 256'hFFFFFFFFFEFFFF7CFDDFFFDE0241FFFFC0003FFA0800300090010FCFDBEB1FFD;
defparam prom_inst_24.INIT_RAM_1F = 256'hFFFFFFFBEFFFFFFE90000FFFFF4003FF961043200000002DFFEF00FD0007FFFF;
defparam prom_inst_24.INIT_RAM_20 = 256'hCE7EF7FFF10300FFFFF0003FFE50031C01000009B7F9980E51881FFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_21 = 256'hFE40000FFFFFFFFFFFFA9000E8000000837FBB80EF19A9FFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_22 = 256'hFFFFFFFDFFFFC031C7800000003FFEC00030057FFFFFFFFFFFFFFFFFFF27F7FF;
defparam prom_inst_24.INIT_RAM_23 = 256'hA3E3FE4002BC0000005FDFFC04003445FFFFFFFFFFFFFFFFFFFD7F4DFEA50880;
defparam prom_inst_24.INIT_RAM_24 = 256'h1101A000009B1FF191000568DFFFFFFFFFFFFFFFFFFFF3F9BFF001003FFFFFFF;
defparam prom_inst_24.INIT_RAM_25 = 256'h00000FBF04002001DBFFFFFFFFFFFFFFFFFFDF2F97D704CA00FFFFFFF231A7FA;
defparam prom_inst_24.INIT_RAM_26 = 256'hBC0080043C3FFFFFFFFFFFFFFFFFFFF93E8FC04101FFFFFFFB0001BFD4060B80;
defparam prom_inst_24.INIT_RAM_27 = 256'h1231FFFFFFFFFFFFFFFFFFFF9EC67C020027FFFFFC01940A3EA0806900000C7F;
defparam prom_inst_24.INIT_RAM_28 = 256'hFFFFFFFFFF85FFFFF9EE85805830DFFFFF8860241DF50121E000005B3FA20010;
defparam prom_inst_24.INIT_RAM_29 = 256'hE9F2FFFFF9C3A65808010FFFFFF9B3FE5C8FA8619FC0001CB9FE200000B03FFF;
defparam prom_inst_24.INIT_RAM_2A = 256'hFF64FFA78140627FFFFF06FFFCA37D48407E000013EDF00472000BFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2B = 256'hF2488006FFFFE6DFFFF3B7EA0963FE4003CFFC140000047FFFFFFFFFFE7FBFDD;
defparam prom_inst_24.INIT_RAM_2C = 256'h1FFFFE4BFFFFD85F50485FF8E21FCF008800008FFFFFFFFFFFDFF7FEFFFF8FFF;
defparam prom_inst_24.INIT_RAM_2D = 256'hBFFFFEC6FA84D03CED3BFFFC200000207FFFFFFFFF1FFF3DFEFFFD3E5B602594;
defparam prom_inst_24.INIT_RAM_2E = 256'h2FD4005FFCE16FFFC00000200FFFFFFFFFF3FF7DFFEFFBF4E77D00293FFFFFD1;
defparam prom_inst_24.INIT_RAM_2F = 256'h1019DAEFF008000018FFFFFFFFFFFFBFFFDFFFFF37B5883112FFFFFC57FFFFF4;
defparam prom_inst_24.INIT_RAM_30 = 256'hF7080200081FFFFFFFFFFFFFDFD9FFFFF35FFC032113FFFFC17FE7FFB0FE2017;
defparam prom_inst_24.INIT_RAM_31 = 256'h0C0B7FFFFFFFFEFFFFFFFFFFC33FBEC0341F7FFFFD07FFFFFD27F30388017FFB;
defparam prom_inst_24.INIT_RAM_32 = 256'hFFFFFFFDFFFFFFFFFC09FF7C0043FFFFFFC2FFF7BFD07FB9B08001BFDD808080;
defparam prom_inst_24.INIT_RAM_33 = 256'hB7FFFFF7FFC03FCF90805FFFFFFD27FFFFFD8FFDDB000007FFFA040000039FFF;
defparam prom_inst_24.INIT_RAM_34 = 256'hFFFE04F9BF258A7FFFFFD07FFFFFD37FE82000003FFE24200C0021FFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_35 = 256'hBCE01C47FFFFFE53FFFFFD27FE660000077FE80004000077FFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_36 = 256'hFFFFFFEC1FFFFF817FF60000001FFE68104000A0BFFFFFFFFFFFFFFC0FFFE035;
defparam prom_inst_24.INIT_RAM_37 = 256'h00FFFFF58FFF23000000BFE0000481203DFFFFFFFFFFFF8A081FFE0054622160;
defparam prom_inst_24.INIT_RAM_38 = 256'h01FFF20000000BFE8400060003FFFFFFFFFFFFFB3803FFF003CFB8171FFFFFFF;
defparam prom_inst_24.INIT_RAM_39 = 256'h000000FFFD000000401FFFFFFFFFFFFFC7C01FFF878CFF0163FFFFFFF56FFFFE;
defparam prom_inst_24.INIT_RAM_3A = 256'hFF6002900009FFFFFFFFFFFFF02C01FFFFFFFDE00FFFFFFFFFB07FFF86DFFE40;
defparam prom_inst_24.INIT_RAM_3B = 256'h00005FFFFFFFFFFFFF0000063FFFFFBF0BDFFFFFFFFD87FFF00BFFF400000009;
defparam prom_inst_24.INIT_RAM_3C = 256'hFFFFFFFFFFF03BC0807FFFFAE9E7FFFFFFFFD1BFFA437FFF680000009FF90000;
defparam prom_inst_24.INIT_RAM_3D = 256'hFFFF879C0C07FFFFCBECFFFFFFFFFE8871002FFFF20000001FFFE00000011AFF;
defparam prom_inst_24.INIT_RAM_3E = 256'h00807FFFFF29FFFFFFFFFFF00C0033FFFFB00000013FFE000020204FFFFFFFFF;
defparam prom_inst_24.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFF5C001CFFBFF90020003FFFE01C000000FFFFFFFFFFFFF879;

pROM prom_inst_25 (
    .DO({prom_inst_25_dout_w[30:0],prom_inst_25_dout[13]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_25.READ_MODE = 1'b1;
defparam prom_inst_25.BIT_WIDTH = 1;
defparam prom_inst_25.RESET_MODE = "SYNC";
defparam prom_inst_25.INIT_RAM_00 = 256'hFFFFFFFFFCE2357FF9FFC800000EFFFF6000011207FFFFFFFFFFFFC6000807FF;
defparam prom_inst_25.INIT_RAM_01 = 256'hFFF22F9FFE0FFE400001FBFFE0003010187FFFFFFFFFFFFA6000007FFFFFFFFF;
defparam prom_inst_25.INIT_RAM_02 = 256'hFF003FF2000C023FFE600000008FFFFFFFFFFFFF9E00300FFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_03 = 256'h900100A7FF80000200007FFFFFFFFFFFFFE00DC0FFFFFFFFFFFFFFFFFFFFC017;
defparam prom_inst_25.INIT_RAM_04 = 256'h1FF98040E0010FFFFFFFFFFFFFF7043C0FFFFFFFFFFFFFFFFFFFFFFFBFE001FF;
defparam prom_inst_25.INIT_RAM_05 = 256'h000003FFFFFFFFFFFFFFC007C1FFFFFFFFFFFFFFFFFFFFFFFFFE200FFCD0E030;
defparam prom_inst_25.INIT_RAM_06 = 256'hFFFFFFFFFFFFF843383FFFFFFFFFFFFFFFFFFFFFFFFFE208FFF3100401FF9000;
defparam prom_inst_25.INIT_RAM_07 = 256'hFFFFFF82A703FFFFFFFFFFFFFFFFFFFFFFFFFE010FFF87A480C7FE200000001F;
defparam prom_inst_25.INIT_RAM_08 = 256'h0AA07FFFFFFFFFFFFFFFFFFFFFFFFFF0007FFF0290103FA000002043FFFFFFFF;
defparam prom_inst_25.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF001FFFF060121BFC100080037FFFFFFFFFFFFFE;
defparam prom_inst_25.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFF801FFFFE50070F9400000200FFFFFFFFFFFFFFF2781FFF;
defparam prom_inst_25.INIT_RAM_0B = 256'hFFFFFFFFF61D01FFFFFA80C23AC00400043FFFFFFFFFFFFFFFF003FFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_0C = 256'hFE03C06FFFFFD022C0E020080002FFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_0D = 256'h9FFFFE80B01E1A381000AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_0E = 256'h00216000400000FFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFF42FE06;
defparam prom_inst_25.INIT_RAM_0F = 256'hC00000DFFFFFFFFFFFFFFFFFFF987FFFFFFFFFFFFFFFFFFFFF17FFFA17FFFFF4;
defparam prom_inst_25.INIT_RAM_10 = 256'h7FFFFFFFFFFFFFFFFFFB3DFFFFFFFFFFFFFFFFFFFC67FFFE019FFFFFA02C2F9C;
defparam prom_inst_25.INIT_RAM_11 = 256'hFFFFFFFFFFFE57CFFFFF61BFFFFFFDFEA0CFFFFFFFFFFFFFFD880868C0304800;
defparam prom_inst_25.INIT_RAM_12 = 256'hFFFFE4B4FFFFE000FFFFFFFC68FFFFFFFFFFFED3FFEC030BA07400001FFFFFFF;
defparam prom_inst_25.INIT_RAM_13 = 256'h4FFFFE0001FFFFF9DFFFFFFFFFFFFFF63FFFE2C21525380041FFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_14 = 256'h001FFFF8DFFFFFFFFFFFFFFF00FFFF00C2F83008040FFFFFFFFFFFFFFFFFFECF;
defparam prom_inst_25.INIT_RAM_15 = 256'h2FFFFFFFFFFFFF48F387FFF83487873A4000FFFFFFFFFFFFFFFFFFEC4DFFFFE0;
defparam prom_inst_25.INIT_RAM_16 = 256'hE00000002F300FFFC810BA0390401FFFFFFFFFFFFFFFFFFE4C9FFFFE0001FFFC;
defparam prom_inst_25.INIT_RAM_17 = 256'hE3E2301FFE0D01FCF4508DBFFFFFFFFFFFFFFFFFFDB3FFFFE0000FFFB7FFFFFF;
defparam prom_inst_25.INIT_RAM_18 = 256'h7FF0090EFF889487FFFFFFFFFFFFFFFFF3E67FFFFE0002FFDBFFFFFF0B040000;
defparam prom_inst_25.INIT_RAM_19 = 256'h77AA2024FFFFFFFFFFFFFFFFFFF14FFFFFE0001FF4FFFFFE11FFFFD998678020;
defparam prom_inst_25.INIT_RAM_1A = 256'h7FFFFFFFFFFFFFFFFFEF39FFFFFE0003F93FFFFFB7FFFFF5D9FFF8412DFF81A4;
defparam prom_inst_25.INIT_RAM_1B = 256'hFFFFFFFFFFFCF73FFFFFE001FE1FFFFFCBFFFFFDFD9AFFE0082FFC3103EF0202;
defparam prom_inst_25.INIT_RAM_1C = 256'hFFFFA267FFFFFF802FC7FFFFF1FFFFFFFCFEC9BFC492FFE0205FF52087FFFFFF;
defparam prom_inst_25.INIT_RAM_1D = 256'hFFFFFFF807E4FFFFF97FFFFFFFFFFFFBFF000FFC3818FF2001BFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_1E = 256'hC17D3FFFFE3FFFFFFFFFFFFFF3E4103FF00817F80014FFFFFFFFFFFFFFFFFFEC;
defparam prom_inst_25.INIT_RAM_1F = 256'hFE2FFFFFFFFFFFFFFFDFB03EFF83443F8000FFFFFFFFFFFFFFFFFFBC9FFFFFFF;
defparam prom_inst_25.INIT_RAM_20 = 256'hFFFFFFFFFFFFFF223FF84105A0000BBFFFFFFFFFFFFFFFE8B3FFFFFFFEDF0FFF;
defparam prom_inst_25.INIT_RAM_21 = 256'hFFFFFFFE17FFC0C10E00007FFFFFFFFFFFFFFFFE1B3FFFFFFFFFE9FFFF97FFFF;
defparam prom_inst_25.INIT_RAM_22 = 256'hF3DFFF00081000097FFFFFFFFFFFFFFF9127FFFFFFFFFD3FFFE1FFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_23 = 256'h0D2180007FFFFFFFFFFFFFFFFF4CFFFFFFFFFFE7FFFDFFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_25.INIT_RAM_24 = 256'h77FFFFFFFFFFFFFFFF4C8FFFFFFFFFF4FFFF3FFFFFFFFFFFFFFFFFFF7FFFFFF0;
defparam prom_inst_25.INIT_RAM_25 = 256'hFFFFFFFFFFE4D9FFFFFFFFFF3FFFDFFFFFFFFFFFFFFFFFFFFFDFFFFF81880400;
defparam prom_inst_25.INIT_RAM_26 = 256'hFFFEC13FFFFFFFFFE3FFFBFFFFFFFFFFFFFFFFFFFFBFFFFFFC05024FE307FFFF;
defparam prom_inst_25.INIT_RAM_27 = 256'hFFFFFFFFFD7FFE7FFFFFFFFFFFFFFFFFFFFCFFFFFFE18003FE703FFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_28 = 256'hFFEFFFC7FFFFFFFFFFFFFFFFFFFFFFBFFFFF0030B7FF85FFFFFFFFFFFFFF8273;
defparam prom_inst_25.INIT_RAM_29 = 256'hFFFFFFFFFFF9FFFFFFFFFEFFFFFFF81F31FFF95FFFFFFFFFFFFFF9E67FFFFFFF;
defparam prom_inst_25.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFF3DFFFFFC28C1DFFE7FFFFFFFFFFFFFFEE4FFFFFFFFFFDFFF9;
defparam prom_inst_25.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFF03E03BFDFFFFFFFFFFFFFFF19CFFFFFFFFFE9FFFBFFFFFFF;
defparam prom_inst_25.INIT_RAM_2C = 256'hFFFFFFFFF02060FFE7FFFFFFFFFFFFFC519FFFFFFFFFEBFFF5FFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_2D = 256'hFFA05847FC1FFFFFFFFFFFFFE693FFFFFFFFFD7FFFBFFFFFFFFFFFC7FFFFFFFF;
defparam prom_inst_25.INIT_RAM_2E = 256'h1FFFFFFFFFFFFFFFF1623FFFFFFFFFAFFFC7FFFFFFFFFFFF7FFFFFFFFFDFFFFF;
defparam prom_inst_25.INIT_RAM_2F = 256'hFFFFFFFFFE04E7FFFFFFFFF5FFFC7FFFFFFFFFFFF7FFFFFFFFFFFFFFFFFD3C18;
defparam prom_inst_25.INIT_RAM_30 = 256'hFF1C8CFFFFFFFFFF5FFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0050BFDFFFF;
defparam prom_inst_25.INIT_RAM_31 = 256'hFFFFFFFFEBFFF5FFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFF41831FCFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_32 = 256'hFE7FFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0182FFFFFFFFFFFFF0323C8F;
defparam prom_inst_25.INIT_RAM_33 = 256'hFFFFFFFFFFFFFC3FFFFFFFFBFFFFFFFFD014C3FFFFFFFFFFFC00CF38FFFFFFFF;
defparam prom_inst_25.INIT_RAM_34 = 256'hFFFFFFF1FFFFFFFFFFFFFFFFFE9C3C3FFFFFFFFFFE001B810FFFFFFFFFC7FFE3;
defparam prom_inst_25.INIT_RAM_35 = 256'h86FFFFFFFFFFFFFFFFF40201FFFFFFFFFFC0036130FFFFFFFFFAFFFE7FFFFFFF;
defparam prom_inst_25.INIT_RAM_36 = 256'hFFFFFFFFFFFFA3910FFFFFFFFFF8003FA20FFFFFFFFFAFFF87FFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_37 = 256'hFFFFFD20816FFFFFFFFF800BE8083FFFFFFFF1FFF8FFFFFFFFFFFFFFFC37FFFF;
defparam prom_inst_25.INIT_RAM_38 = 256'h1643FFFFFFFFF800B78043FFFFFFFF5FFF1FFFFFFFFFFFFFFFF02FFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_39 = 256'hFFFFFF0097B8003FFFFFFFE3FFF1FFFFFFFFFFFFFFFF8715FFFFFFFFFFFFFFE8;
defparam prom_inst_25.INIT_RAM_3A = 256'h210F0011FFFFFFFF3FFE3FFFFFFFFFFFFFFFFE017BFD5FFFFFFFFFFF4A591FFF;
defparam prom_inst_25.INIT_RAM_3B = 256'h9FFFFFFFCFFFE3FFFFFFFFFFFFFFCFF000180FFFFFFFFFFFFA0500FFFFFFFFF0;
defparam prom_inst_25.INIT_RAM_3C = 256'hFF7FFC7FFFFFFFFFFFFFFC1FF8000FFFFFFFFFFFFFD148C7FFFFFFFF0241E803;
defparam prom_inst_25.INIT_RAM_3D = 256'hFFFFFFFFFFFFFD803FF8CFFFFFFFFFFFFFFE92201FFFFFFFC000740039FFFFFF;
defparam prom_inst_25.INIT_RAM_3E = 256'hFFFFFE4000FFFFFFFFFFFFFFFFFFF41383FFFFFFFE84A4C8019FFFFFFFDFFFC7;
defparam prom_inst_25.INIT_RAM_3F = 256'h0003FFFFFFFFFFFFFFFFFFA4C01FFFFFFFAC43780059FFFFFFF8FFFC7FFFFFFF;

pROM prom_inst_26 (
    .DO({prom_inst_26_dout_w[30:0],prom_inst_26_dout[14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_26.READ_MODE = 1'b1;
defparam prom_inst_26.BIT_WIDTH = 1;
defparam prom_inst_26.RESET_MODE = "SYNC";
defparam prom_inst_26.INIT_RAM_00 = 256'h000000000008FFFFFDFFFFFFC4000000000020C2002201208000000000000001;
defparam prom_inst_26.INIT_RAM_01 = 256'h000DFFFFFEDFFFFFE79800000500000200204000000000000000000000000000;
defparam prom_inst_26.INIT_RAM_02 = 256'hFFE1FFFFFFE6A0400000033B9FB5FC2124000000000000000000000000000000;
defparam prom_inst_26.INIT_RAM_03 = 256'hFFFFFA001860109BEFFC57925650000000000000000000000000000000001FFF;
defparam prom_inst_26.INIT_RAM_04 = 256'h13A8127E7FFFF7EB94BE000000000000000000000000000000000DFFFFE907FF;
defparam prom_inst_26.INIT_RAM_05 = 256'hFDFDEFFDB2DF3A00000000000000000000000000000005FFFFFF000FFFFFFFA3;
defparam prom_inst_26.INIT_RAM_06 = 256'hF265C5080000000000000000000000000000017BFFFF00001DFFFFCF380FE2EF;
defparam prom_inst_26.INIT_RAM_07 = 256'h1800000000000000000000000000000BF7FFFA0000FFFFFFFFC7B9DFFFFFDFFF;
defparam prom_inst_26.INIT_RAM_08 = 256'h0000000000000000000000019FFFFE180201FFFFEAC037FF1FFFFFFFFFDC39E0;
defparam prom_inst_26.INIT_RAM_09 = 256'h00000000000000016FFFFF40A04007FF3FA2039FFFFFFFFFFFFEF40C9A000000;
defparam prom_inst_26.INIT_RAM_0A = 256'h0000000007FFFF5002900037FA7AC017FFFFFBEFFEFF6F3C6640000000000000;
defparam prom_inst_26.INIT_RAM_0B = 256'h007BFFE8000C0000FCA60C013FFFFFDFFFFFFFEAA60400000000000000000000;
defparam prom_inst_26.INIT_RAM_0C = 256'h800088002000104041FFFFF9BFFDFFFFFC6C4000010000000000000000000002;
defparam prom_inst_26.INIT_RAM_0D = 256'h0C078000001BFFFFDF339FDFFF7F002300000000000000000000000000003FFF;
defparam prom_inst_26.INIT_RAM_0E = 256'h0001FFFFFBFEFFDFFFF0602000000080000000000000000000004FFFE0002460;
defparam prom_inst_26.INIT_RAM_0F = 256'hFFFFFDEFFFFF4E00400000000000000000000000000000DFF800080080001000;
defparam prom_inst_26.INIT_RAM_10 = 256'hF77FFD90C0400100000000000000000000000017FF0081000340004000001FFF;
defparam prom_inst_26.INIT_RAM_11 = 256'h884000008000000000000000000000113F40004000100000000001FFFFE003BF;
defparam prom_inst_26.INIT_RAM_12 = 256'h0000000000000000000000000EF80000800030008000003FFFF43FB7FFFFFFC2;
defparam prom_inst_26.INIT_RAM_13 = 256'h000000000000000000FA00002000014020000001FFFF1FE43F7FCFEF40040000;
defparam prom_inst_26.INIT_RAM_14 = 256'h000000000009800040801212048000003FFFC7ADE3FFFEFFBE40800600000000;
defparam prom_inst_26.INIT_RAM_15 = 256'h0000F900102602000800000007FF79FF8017FFFFFFF014000203240000000000;
defparam prom_inst_26.INIT_RAM_16 = 256'h0400A89001140000007FFF1F0E60FFFFFFFF8880212440000000000000000000;
defparam prom_inst_26.INIT_RAM_17 = 256'h00108000003FFFF0E06007FFFFFFF9200A009800000000000000000000001E81;
defparam prom_inst_26.INIT_RAM_18 = 256'h00017FEE0788000FFFFFFDE0000010C100000000000000000000001010500221;
defparam prom_inst_26.INIT_RAM_19 = 256'hE03A00103FFFFFDF000009A52100000000000000000000400040000800008000;
defparam prom_inst_26.INIT_RAM_1A = 256'h03FFE3FFF7004011024000000000000000000000D00000000200248000001FFF;
defparam prom_inst_26.INIT_RAM_1B = 256'hBFFB00A11040000000000000000000000080480021080408000002FFFC01C01C;
defparam prom_inst_26.INIT_RAM_1C = 256'h00342C3DF00000000000000000010010000260208000003FFFF0080EE03FFF0B;
defparam prom_inst_26.INIT_RAM_1D = 256'h7F40000000000000000E0004810008A009100003FFFF80036540FFC7DDC7D420;
defparam prom_inst_26.INIT_RAM_1E = 256'h000000000100000212200020000900003FFFC00048404FFF6FFEF0302414E002;
defparam prom_inst_26.INIT_RAM_1F = 256'h00000002084000010000100000BFFC00021340DFFFFFFFD20010FF02FFF80000;
defparam prom_inst_26.INIT_RAM_20 = 256'h0800080000010100000FFFC000704303FEFFFFF6480667F1AE77E00000000000;
defparam prom_inst_26.INIT_RAM_21 = 256'h0150001000000000000390C017FFFFFF7C80447F10E656000000000000000000;
defparam prom_inst_26.INIT_RAM_22 = 256'h0000000008000C33C07FFFFFFFC0013FFFCFFA80000000000000000004300000;
defparam prom_inst_26.INIT_RAM_23 = 256'h884000608283FFFFFFA02003FBFFCBBA00000000000000000000409201050081;
defparam prom_inst_26.INIT_RAM_24 = 256'h11005FFFFF64E00E6EFFFA972000000000000000000002004000410000000000;
defparam prom_inst_26.INIT_RAM_25 = 256'hFFFFF040FBFFDFFE240000000000000000000080012800080400000000001803;
defparam prom_inst_26.INIT_RAM_26 = 256'h43FF7FFBC3C0000000000000000000000504000000D00000000000001C26847F;
defparam prom_inst_26.INIT_RAM_27 = 256'hEDCE0000000000000000000000000402000900000100E80040E0A016FFFFF380;
defparam prom_inst_26.INIT_RAM_28 = 256'h00000000004A000045140100081410000000E038000700A01FFFFFA4C05DFFEF;
defparam prom_inst_26.INIT_RAM_29 = 256'h0A02C00001000800000101000004100060203861903FFFE34601DFFFFF4FC000;
defparam prom_inst_26.INIT_RAM_2A = 256'h00840000014800100000020000C001C82001FFFFEC120FFB8DFFF40000000000;
defparam prom_inst_26.INIT_RAM_2B = 256'h00008400000000400002000E196001BFFC3003EBFFFFFB80000000000260BC3E;
defparam prom_inst_26.INIT_RAM_2C = 256'h4000000000001000705840071DE030FF77FFFF7000000000001F0FC2E0000801;
defparam prom_inst_26.INIT_RAM_2D = 256'h800000800384902212C40003DFFFFFDF8000000000E3F0FE3E00024004282080;
defparam prom_inst_26.INIT_RAM_2E = 256'h001C1060011E90003FFFFFDFF000000000131F8383E000111009420848000010;
defparam prom_inst_26.INIT_RAM_2F = 256'h000025100FF7FFFFE70000000001F0381C1C0000604000150400000000000006;
defparam prom_inst_26.INIT_RAM_30 = 256'h08F7FDFFF7E0000000001FC3E1E1800100040001000000000000180020006018;
defparam prom_inst_26.INIT_RAM_31 = 256'hF3F48000000000FF1FFFF8000480000010080000001000000100030206000004;
defparam prom_inst_26.INIT_RAM_32 = 256'h00000003FFFFFF8000120000040100000010800840100039C3000040227F7F7F;
defparam prom_inst_26.INIT_RAM_33 = 256'h4FFFFFF00000200000B400000001080000010801E00000000005FBFFFFFC6000;
defparam prom_inst_26.INIT_RAM_34 = 256'h000001010500C00000001040000010800F0000000001DBDFF3FFDE0000000000;
defparam prom_inst_26.INIT_RAM_35 = 256'h45040D00000000800000000800500000008017FFFBFFFF8800000000003FFFFF;
defparam prom_inst_26.INIT_RAM_36 = 256'h00000008000000000007000000000197EFBFFF5F400000000000FFFFFC000000;
defparam prom_inst_26.INIT_RAM_37 = 256'h41000000200030000000401FFFFB7EDFC2000000000007FFF040000000042060;
defparam prom_inst_26.INIT_RAM_38 = 256'h00000300000010017BFFF9FFFC00000000000000FF0000000080040400000000;
defparam prom_inst_26.INIT_RAM_39 = 256'h0000000002FFFFFFBFE00000000000000FE00000000000000000000006000000;
defparam prom_inst_26.INIT_RAM_3A = 256'h009FFD6FFFF60000000000000010008000000800200000000020000000400070;
defparam prom_inst_26.INIT_RAM_3B = 256'hFFFFA00000000000008000080000000104000000000104001008000700000000;
defparam prom_inst_26.INIT_RAM_3C = 256'h000000000000000040000000148000000000180008010000700000000006FFFF;
defparam prom_inst_26.INIT_RAM_3D = 256'h000000000000000000400000000000820800E0000300000000001FFFFFFEE500;
defparam prom_inst_26.INIT_RAM_3E = 256'h0040000000000000000000040000100000380000000001FFFFDFDFB000000000;
defparam prom_inst_26.INIT_RAM_3F = 256'h000000000000000060010C004001C0000000001FE3FFFFFF0000000000000800;

pROM prom_inst_27 (
    .DO({prom_inst_27_dout_w[30:0],prom_inst_27_dout[14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_27.READ_MODE = 1'b1;
defparam prom_inst_27.BIT_WIDTH = 1;
defparam prom_inst_27.RESET_MODE = "SYNC";
defparam prom_inst_27.INIT_RAM_00 = 256'h0000000000C01B0006000E00000140009FFFFEEDF80000000000000000080000;
defparam prom_inst_27.INIT_RAM_01 = 256'h0003F38001F00070000000001FFFCFEFE7800000000000040001000000000000;
defparam prom_inst_27.INIT_RAM_02 = 256'h00FFC00380000000019FFFFFFF70000000000000200010000000000000000000;
defparam prom_inst_27.INIT_RAM_03 = 256'h1C00006C007FFFFDFFFF80000000000000000FC0000000000000000000000010;
defparam prom_inst_27.INIT_RAM_04 = 256'h00067FBF1FFEF0000000000000000C3C000000000000000000000000001FFE00;
defparam prom_inst_27.INIT_RAM_05 = 256'hFFFFFC000000000000000805C000000000000000000000000001DFF000E00010;
defparam prom_inst_27.INIT_RAM_06 = 256'h00000000000000C218000000000000000000000000001DF70003E00C01006FFF;
defparam prom_inst_27.INIT_RAM_07 = 256'h00000003030000000000000000000000000001FEF00007C880C001DFFFFFFFE0;
defparam prom_inst_27.INIT_RAM_08 = 256'h0DE0000000000000000000000000000FFF8000035030005FFFFFDFBC00000000;
defparam prom_inst_27.INIT_RAM_09 = 256'h0000000000000000000000000FFE00000A0A20403EFFF7FFC800000000000000;
defparam prom_inst_27.INIT_RAM_0A = 256'h0000000000000000007FE00000720F006BFFFFFDFF0000000000000000780000;
defparam prom_inst_27.INIT_RAM_0B = 256'h000000000402FE0000038202453FFBFFFBC00000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0C = 256'h02003F90000018A2C31FDFF7FFFD000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0D = 256'h600000C08081E5C7EFFF50000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0E = 256'h28309FFFBFFFFF000000000000000000004000000000000000000000002601F9;
defparam prom_inst_27.INIT_RAM_0F = 256'h3FFFFF20000000000000000000508000000000000000000002300005E8000006;
defparam prom_inst_27.INIT_RAM_10 = 256'h800000000000000000072000000000000000000008200001FE60000030202063;
defparam prom_inst_27.INIT_RAM_11 = 256'h00000000000006000000004000000200C1C0000000000000018A0C173FCFB7FF;
defparam prom_inst_27.INIT_RAM_12 = 256'h000006800000100000000004180000000000012C000C00085F8BFFFFE0000000;
defparam prom_inst_27.INIT_RAM_13 = 256'hC0000000020000044000000000000009C00062430ADAC7FFBE00000000000000;
defparam prom_inst_27.INIT_RAM_14 = 256'h001000004000000000000000FF0003000207CFF7FBF0000000000000000002D8;
defparam prom_inst_27.INIT_RAM_15 = 256'h60000000000000700C78001814C078C5BFFF0000000000000000001A8C000000;
defparam prom_inst_27.INIT_RAM_16 = 256'h3000000010CFF000C82085FC6FBFE00000000000000000019580000000000000;
defparam prom_inst_27.INIT_RAM_17 = 256'hE01DCFE0060410030BAF72400000000000000000461000000000100010000000;
defparam prom_inst_27.INIT_RAM_18 = 256'h80320D0100776B78000000000000000006020000000000004800000107000000;
defparam prom_inst_27.INIT_RAM_19 = 256'h0855DFDB0000000000000000000CC00000200020040000013000000000007FDF;
defparam prom_inst_27.INIT_RAM_1A = 256'h800000000000000000109800000000040100000010000000000007BED20183A4;
defparam prom_inst_27.INIT_RAM_1B = 256'h00000000000003000000100080000000480000000000001FF7D00CB14010FDFD;
defparam prom_inst_27.INIT_RAM_1C = 256'h00000060000000000000000004000000000000003B6D006028400ADF78000000;
defparam prom_inst_27.INIT_RAM_1D = 256'h0000000800040000090000000000000000FFF0003C0800DFFE40000000000000;
defparam prom_inst_27.INIT_RAM_1E = 256'h000000000080000000000000000BEFC0100A1007FFEB0000000000000000000C;
defparam prom_inst_27.INIT_RAM_1F = 256'h002000000000000000004FC1008242007FFF0000000000000000000180000000;
defparam prom_inst_27.INIT_RAM_20 = 256'h00000000000000DDC00040845FFFF44000000000000000141000000000000000;
defparam prom_inst_27.INIT_RAM_21 = 256'h00000001E800008981FFFF800000000000000002030000000000100000400000;
defparam prom_inst_27.INIT_RAM_22 = 256'h0C200110682FFFF6800000000000000000600000000002000014000000000000;
defparam prom_inst_27.INIT_RAM_23 = 256'h1D207FFF80000000000000000024000000000040000100000000000000000000;
defparam prom_inst_27.INIT_RAM_24 = 256'h8800000000000000002080000000000000014000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_25 = 256'h00000000001018000000000000000000000000000000000000200000058A0BFF;
defparam prom_inst_27.INIT_RAM_26 = 256'h00020B000000000000000200000000000000000000000000000542301CF80000;
defparam prom_inst_27.INIT_RAM_27 = 256'h00000000010000400000000000000000000000000001E0C0018FC00000000000;
defparam prom_inst_27.INIT_RAM_28 = 256'h0000000000000000000000000000004000000000A8007A000000000000000130;
defparam prom_inst_27.INIT_RAM_29 = 256'h00000000000000000000000000000017210006A0000000000000000600000000;
defparam prom_inst_27.INIT_RAM_2A = 256'h000000000000000020000002801A00180000000000000000C000000000080001;
defparam prom_inst_27.INIT_RAM_2B = 256'h000000000000000101A4040200000000000000004C0000000000000020000000;
defparam prom_inst_27.INIT_RAM_2C = 256'h0000000000A16100180000000000000289800000000008000400000000000000;
defparam prom_inst_27.INIT_RAM_2D = 256'h0020404803E00000000000004130000000000100000000000000000000000000;
defparam prom_inst_27.INIT_RAM_2E = 256'h6000000000000000009600000000004000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_2F = 256'h0000000000226000000000000000000000000000000000000000000000013810;
defparam prom_inst_27.INIT_RAM_30 = 256'h00004C0000000000400020000000000000000000000000000000000108020000;
defparam prom_inst_27.INIT_RAM_31 = 256'h000000001000080000000000000000000000000000000040A100300000000000;
defparam prom_inst_27.INIT_RAM_32 = 256'h0000000000000000000000000000000000000002414200000000000010300180;
defparam prom_inst_27.INIT_RAM_33 = 256'h000000000000000000000000000000001078C000000000000400809800000000;
defparam prom_inst_27.INIT_RAM_34 = 256'h000000000000000000000000009E382000000000000010130000000000100000;
defparam prom_inst_27.INIT_RAM_35 = 256'h0000000000000000000402850000000000000203F00000000000000100000000;
defparam prom_inst_27.INIT_RAM_36 = 256'h0000000000002350880000000000000062000000000020000000000000000000;
defparam prom_inst_27.INIT_RAM_37 = 256'h00000120A15000000000000C1408000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_38 = 256'h2462000000000803000040000000004000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_39 = 256'h00000000E0480200000000000000000000000000000000000000000000000008;
defparam prom_inst_27.INIT_RAM_3A = 256'h3E0000300000000080000000000000000000000000000000000000004F5B1000;
defparam prom_inst_27.INIT_RAM_3B = 256'h8000000008000000000000000000400000000000000000000205428000000010;
defparam prom_inst_27.INIT_RAM_3C = 256'h020000000000000000000C000000000000000000001128040000000103801802;
defparam prom_inst_27.INIT_RAM_3D = 256'h0000000000000580000000000000000000009210200000000038038028000000;
defparam prom_inst_27.INIT_RAM_3E = 256'h0000006000000000000000000000041A82000000028700380280000000100000;
defparam prom_inst_27.INIT_RAM_3F = 256'h0000000000000000000000264000000000307807004800000000000000000000;

pROM prom_inst_28 (
    .DO({prom_inst_28_dout_w[30:0],prom_inst_28_dout[15]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_28.READ_MODE = 1'b1;
defparam prom_inst_28.BIT_WIDTH = 1;
defparam prom_inst_28.RESET_MODE = "SYNC";
defparam prom_inst_28.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_28.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC07FFFFFFFFF;
defparam prom_inst_28.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFE003FFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFF8121FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFE1FFFFFFFFFE007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_16 = 256'hFFFFFFFFFFF81FFFFFFFFFE0F181FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_17 = 256'hFFFF01FFFFFFFFFF1F800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_18 = 256'hFFFFFFFFF870007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFF;
defparam prom_inst_28.INIT_RAM_19 = 256'hFFC40007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFF01F;
defparam prom_inst_28.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFFFFFFF901FFFFFFFF;
defparam prom_inst_28.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FFFFFFFFF103FFFFFFFFFFE0003;
defparam prom_inst_28.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FFFFFFFFC107FFFFFFFFFFF0001FFFFFFF;
defparam prom_inst_28.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFF033FFFFFFF810CFFFFFFFFFFF809ABFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1E = 256'hFFFFFFFFFFFFFF810FFFFFFF01B0FFFFFFFFFFFC37BFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1F = 256'hFFFFFFFC103FFFFFE01E0FFFFFFFFFFFE1ECBFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_20 = 256'hB181FFFFFE00C0FFFFFFFFFFFF8FBCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_21 = 256'hFE20380FFFFFFFFFFFFC6F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_22 = 256'hFFFFFFFFC7FFF3CC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8C80FFF;
defparam prom_inst_28.INIT_RAM_23 = 256'h0007FF9F7D7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3806FFFC20700;
defparam prom_inst_28.INIT_RAM_24 = 256'hEE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0C063FF830D81FFFFFFF;
defparam prom_inst_28.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07060FE033183FFFFFF800027FC;
defparam prom_inst_28.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE06C203C03E180FFFFFF000003FE3D97FFF;
defparam prom_inst_28.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFF063301801C190FFFFFE0000003F1F5FFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFF820B00C0300A0FFFFFC01FC003F8FE5FFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_29 = 256'hF7FD3FFFF630700C0700C0FFFFF80FFF801FC79E6FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2A = 256'hFF1B01C0C0B0180FFFFF81FFFF007E379FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2B = 256'h0C330381FFFFF03FFFFC07F1E69FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD9F43E3;
defparam prom_inst_28.INIT_RAM_2C = 256'h3FFFFF07FFFFE01F8FA7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0F03D1FF8701E;
defparam prom_inst_28.INIT_RAM_2D = 256'h7FFFFF00FC7B2FC1FFFFFFFFFFFFFFFFFFFFFFFFFFFC0F83C1FF8181B8C61848;
defparam prom_inst_28.INIT_RAM_2E = 256'h0FE3EF8000FFFFFFFFFFFFFFFFFFFFFFFFECE0FE7C1FFC0E08E6819087FFFFE0;
defparam prom_inst_28.INIT_RAM_2F = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFE0FC7E3E3FFC09883F00A09FFFFFE0FFFFFF8;
defparam prom_inst_28.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFE03C1E1E7FFE0CE80E00C0FFFFFFE0FFFFFFC0FF9FE0;
defparam prom_inst_28.INIT_RAM_31 = 256'hFFFFFFFFFFFFFF00E00007FFF843C0600807FFFFFE0FFFFFFE07FCFC00000FFF;
defparam prom_inst_28.INIT_RAM_32 = 256'hFFFFFFFE0000007FFFE40C060380FFFFFFE07FFFFFE07FC60000003FFFFFFFFF;
defparam prom_inst_28.INIT_RAM_33 = 256'hF800000FFFFFC07060483FFFFFFE07FFFFFE07FE00000001FFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_34 = 256'hFFFFFE06C21807FFFFFFE03FFFFFE07FF00000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_35 = 256'h223300FFFFFFFF03FFFFFE07FF800000007FFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam prom_inst_28.INIT_RAM_36 = 256'hFFFFFFF03FFFFFC0FFF800000007FFFFFFFFFFFFFFFFFFFFFFFF000003FFFFF8;
defparam prom_inst_28.INIT_RAM_37 = 256'h80FFFFF81FFFC00000003FFFFFFFFFFFFFFFFFFFFFFFF800003FFFFFE31BC09F;
defparam prom_inst_28.INIT_RAM_38 = 256'h03FFFC00000003FFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFF30780BFFFFFFFF;
defparam prom_inst_28.INIT_RAM_39 = 256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFF80000FFFFFFF0180FFFFFFFFF80FFFFF;
defparam prom_inst_28.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFF0181FFFFFFFFFC0FFFFE03FFF80;
defparam prom_inst_28.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF000007FFFFFFC083FFFFFFFFFE03FFE007FFF800000003;
defparam prom_inst_28.INIT_RAM_3C = 256'hFFFFFFFFFFF000003FFFFFFF087FFFFFFFFFE03FF000FFFF800000003FFFFFFF;
defparam prom_inst_28.INIT_RAM_3D = 256'hFFFF000003FFFFFFFC9FFFFFFFFFFF0032001FFFFC00000003FFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_3E = 256'h003FFFFFFFFFFFFFFFFFFFF800000FFFFFC00000003FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFF800003FFFFFE00000003FFFFFFFFFFFFFFFFFFFFFFFFF000;

pROM prom_inst_29 (
    .DO({prom_inst_29_dout_w[30:0],prom_inst_29_dout[15]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_29.READ_MODE = 1'b1;
defparam prom_inst_29.BIT_WIDTH = 1;
defparam prom_inst_29.RESET_MODE = "SYNC";
defparam prom_inst_29.INIT_RAM_00 = 256'hFFFFFFFFFF0000FFFFFFF00000003FFFFFFFFFFFFFFFFFFFFFFFFF800007FFFF;
defparam prom_inst_29.INIT_RAM_01 = 256'hFFFC007FFFFFFF80000007FFFFFFFFFFFFFFFFFFFFFFFFF80000FFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_02 = 256'hFFFFFFFC0000007FFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_03 = 256'hE0000013FFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_29.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF803C3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFF7F83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000F;
defparam prom_inst_29.INIT_RAM_06 = 256'hFFFFFFFFFFFFFF3C07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FEFFFFFF;
defparam prom_inst_29.INIT_RAM_07 = 256'hFFFFFFFC00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007F3FFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_08 = 256'hF01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FCFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F4DFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF8DF0FFFFFFFFFFFFFFFFFFFFFFFFFFFF87FFFF;
defparam prom_inst_29.INIT_RAM_0B = 256'hFFFFFFFFF81FFFFFFFFC7D3DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_0C = 256'hFC01FFFFFFFFE75D3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_0D = 256'hFFFFFF3F4F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_0E = 256'hD7CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFE01FFFF;
defparam prom_inst_29.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFC0FFFFFFFFFFFF9;
defparam prom_inst_29.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFF803FFFFFFFFFFFFFFFFFFF01FFFFFFFFFFFFFCFD3DFFF;
defparam prom_inst_29.INIT_RAM_11 = 256'hFFFFFFFFFFFF203FFFFF803FFFFFFFFF003FFFFFFFFFFFFFFE75F3FFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_12 = 256'hFFFFF043FFFFE0007FFFFFF807FFFFFFFFFFFFFFFFF3FCF7FFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_13 = 256'h3FFFFE0001FFFFF83FFFFFFFFFFFFFFFFFFF9D3CFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_14 = 256'h000FFFFC3FFFFFFFFFFFFFFFFFFFFCFF3DFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_29.INIT_RAM_15 = 256'h1FFFFFFFFFFFFF80FFFFFFE7CB3FFFFFFFFFFFFFFFFFFFFFFFFFFFC103FFFFC0;
defparam prom_inst_29.INIT_RAM_16 = 256'hC00000000FFFFFFF37CF7FFFFFFFFFFFFFFFFFFFFFFFFFFC207FFFFC0000FFFE;
defparam prom_inst_29.INIT_RAM_17 = 256'h1FFFFFFFF9F2EFFFFFFFFFFFFFFFFFFFFFFFFFFF800FFFFFC0000FFF0FFFFFFF;
defparam prom_inst_29.INIT_RAM_18 = 256'hFFCDF2FFFFFFFFFFFFFFFFFFFFFFFFFFF801FFFFFC0001FF87FFFFFE00FFFFFF;
defparam prom_inst_29.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF003FFFFFC0001FE3FFFFFE0FFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFE007FFFFFE0003F8FFFFFF0FFFFFFFFFFFFFFFFFFE7C1B;
defparam prom_inst_29.INIT_RAM_1B = 256'hFFFFFFFFFFFE00FFFFFFE0007E7FFFFF87FFFFFFFFFFFFFFFFFFF34EBFFFFFFF;
defparam prom_inst_29.INIT_RAM_1C = 256'hFFFFC01FFFFFFF001F9FFFFFE3FFFFFFFFFFFFFFFFFFFF9FC7BFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_1D = 256'hFFFFFFF003F3FFFFF0FFFFFFFFFFFFFFFFFFFFFFC3E7FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_1E = 256'h80FCFFFFFC7FFFFFFFFFFFFFFFFFFFFFEFF1EFFFFFFFFFFFFFFFFFFFFFFFF803;
defparam prom_inst_29.INIT_RAM_1F = 256'hFF1FFFFFFFFFFFFFFFFFFFFFFF7CB9FFFFFFFFFFFFFFFFFFFFFFFF007FFFFFFF;
defparam prom_inst_29.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFBE7BFFFFFFFFFFFFFFFFFFFFFFE00FFFFFFFFC3FBFFF;
defparam prom_inst_29.INIT_RAM_21 = 256'hFFFFFFFFFFFFFF367FFFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFFE7FFFF8FFFFF;
defparam prom_inst_29.INIT_RAM_22 = 256'hFFFFFEEF97FFFFFFFFFFFFFFFFFFFFFFC01FFFFFFFFFFCFFFFE3FFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_23 = 256'hE0DFFFFFFFFFFFFFFFFFFFFFF803FFFFFFFFFF9FFFF8FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFF007FFFFFFFFFFBFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_25 = 256'hFFFFFFFFFFE007FFFFFFFFFF7FFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFA75FFFF;
defparam prom_inst_29.INIT_RAM_26 = 256'hFFFC00FFFFFFFFFFEFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFA3DFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_27 = 256'hFFFFFFFFFCFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFE1F3FFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_28 = 256'hFF9FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF5FFFFFFFFFFFFFFFFFFFC00F;
defparam prom_inst_29.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0CEFFFFFFFFFFFFFFFFFFF801FFFFFFFF;
defparam prom_inst_29.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFD73E7FFFFFFFFFFFFFFFFFF003FFFFFFFFFF3FFFC;
defparam prom_inst_29.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFEFC1BFFFFFFFFFFFFFFFFFFE003FFFFFFFFFF7FFF9FFFFFFF;
defparam prom_inst_29.INIT_RAM_2C = 256'hFFFFFFFFFF5E9FFFFFFFFFFFFFFFFFFC007FFFFFFFFFE7FFF3FFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2D = 256'hFFDFA7BFFFFFFFFFFFFFFFFF800FFFFFFFFFFCFFFE7FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFF801FFFFFFFFFF9FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2F = 256'hFFFFFFFFFF001FFFFFFFFFFBFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC3E7;
defparam prom_inst_29.INIT_RAM_30 = 256'hFFE003FFFFFFFFFF3FFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F7FFFFFF;
defparam prom_inst_29.INIT_RAM_31 = 256'hFFFFFFFFE7FFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBE5CFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_32 = 256'hFEFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDBE3DFFFFFFFFFFFFEFCC007F;
defparam prom_inst_29.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF833FFFFFFFFFFFFBFF0007FFFFFFFF;
defparam prom_inst_29.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF61C3DFFFFFFFFFFFFFE000FFFFFFFFFFCFFFEF;
defparam prom_inst_29.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFBFC7AFFFFFFFFFFFFFC000FFFFFFFFFFDFFFCFFFFFFFF;
defparam prom_inst_29.INIT_RAM_36 = 256'hFFFFFFFFFFFFDC2E77FFFFFFFFFFFFC01DFFFFFFFFFF9FFFDFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_37 = 256'hFFFFFEDF1EBFFFFFFFFFFFF003F7FFFFFFFFFBFFFBFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_38 = 256'hC99DFFFFFFFFF7FC007FBFFFFFFFFF3FFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_39 = 256'hFFFFFFFF0007FDFFFFFFFFF7FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;
defparam prom_inst_29.INIT_RAM_3A = 256'hC000FFCFFFFFFFFE7FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB0A4EFFF;
defparam prom_inst_29.INIT_RAM_3B = 256'h7FFFFFFFE7FFEFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFDFA3D7FFFFFFFEF;
defparam prom_inst_29.INIT_RAM_3C = 256'hFCFFFEFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFEE973BFFFFFFFEFC0007FC;
defparam prom_inst_29.INIT_RAM_3D = 256'hFFFFFFFFFFFFFA7FFFFFFFFFFFFFFFFFFFFF6DCFFFFFFFFFFFC0007FC7FFFFFF;
defparam prom_inst_29.INIT_RAM_3E = 256'hFFFFFF9FFFFFFFFFFFFFFFFFFFFFFBE47DFFFFFFFD780007FC7FFFFFFFCFFFDF;
defparam prom_inst_29.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFD93FFFFFFFFFC38000FF87FFFFFFFDFFFDFFFFFFFF;

pROMX9 promx9_inst_30 (
    .DO({promx9_inst_30_dout_w[26:0],promx9_inst_30_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_35),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_30.READ_MODE = 1'b1;
defparam promx9_inst_30.BIT_WIDTH = 9;
defparam promx9_inst_30.RESET_MODE = "SYNC";
defparam promx9_inst_30.INIT_RAM_00 = 288'hCAE572B95CAE56EB95BADD6EB75BADD6EB75AAD56AB54AA4D269138A2CE9305D1B81C922;
defparam promx9_inst_30.INIT_RAM_01 = 288'h9A349C6D289CD2AB54BADD6EB75CAE572B95CAE572B95BAE572B95CAE572B95CAE572B95;
defparam promx9_inst_30.INIT_RAM_02 = 288'hCAE572B95CAE572B95CAE572B95CADD72B75BA1C21313BADD6EB75BADD6EB75BADD6AB54;
defparam promx9_inst_30.INIT_RAM_03 = 288'hE350F0BE452A994AA663319CCC62359144EBE7245E734AA556EB75BADD72B95CAE572B95;
defparam promx9_inst_30.INIT_RAM_04 = 288'hDB6DB6DB6DB6DB6D96CADD2EAD223A9AD8EAF3384CA4532A1A0784D2B0A08E371D1608C2;
defparam promx9_inst_30.INIT_RAM_05 = 288'h724924B2482C160B2592C964B2592C9A8D95DAE576D95DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_06 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6CACD31B04;
defparam promx9_inst_30.INIT_RAM_07 = 288'hCAED76B95DAEDB2D96DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB75B6DB6;
defparam promx9_inst_30.INIT_RAM_08 = 288'h5140A46C2B248E47228140A44E29140A06E27161140E5A9DDAEB95BAE56EB75CAE572B95;
defparam promx9_inst_30.INIT_RAM_09 = 288'hCAE572B95CAE572B95CAE56EB95BAE56EB75BADD6EB75AA552AB348A451E6D36949F0803;
defparam promx9_inst_30.INIT_RAM_0A = 288'hBAD56A9549A79D12D29A552AB54BADD6EB75CADD72B95CAE572B95CAE572B95CAE572B95;
defparam promx9_inst_30.INIT_RAM_0B = 288'hCAE572B95CAE572B95CAE572B95CAE572B95BAE56EB75AA21ED934BADD6EB75BADD6EB75;
defparam promx9_inst_30.INIT_RAM_0C = 288'h91B8F4D84B1E1786A6532994CC67339DCE45F2A8B8F6D182CA2734AADD6EB75CAE572B95;
defparam promx9_inst_30.INIT_RAM_0D = 288'hDB6DB6DB6DB6DB6D95DAE572B95BA9C14EC7C4E241CA7331948A6532997CB64B25138D03;
defparam promx9_inst_30.INIT_RAM_0E = 288'hDB656278E92C124B2582C964B25A2C964B2592C974FB5DB6576DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_0F = 288'hDB75BADD6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6EB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_10 = 288'hCAE572B95CAE572B95DAEDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_11 = 288'h6378C848380D0E4783C238AC923A1C8A05438140A050260A8585845149EE975BADD6EB95;
defparam promx9_inst_30.INIT_RAM_12 = 288'hCAE572B95CAE572B95CAE572B75BAE56EB75BADD6EB75BAD56AB54AA4D268F389BCDA492;
defparam promx9_inst_30.INIT_RAM_13 = 288'hBADD6EB75BAD56A95489B0CE2F39A552AB54BADD6EB75CAE572B95CAE572B95CAE572B95;
defparam promx9_inst_30.INIT_RAM_14 = 288'hCAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE56EB759A3205F54BADD6EB75;
defparam promx9_inst_30.INIT_RAM_15 = 288'h81D130B2381D128965A22194CA6632994CE773B9C49A350A8E17EF48BCE6954AADD6EB75;
defparam promx9_inst_30.INIT_RAM_16 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6D95CAE56EBAD443A45E7027A181AA542A194CA5429950DE5;
defparam promx9_inst_30.INIT_RAM_17 = 288'hDB6DB6DB6DB6DAEB5407D15C925A2C164B2592C964B2592C9A2995CAE576DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_18 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DAEDB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_19 = 288'hBADD32B95CAE572B95CAE572B95CAE576BB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_1A = 288'h79B4924C532F090302B1E130984C261182C2B240A05028140A05028138542807168D07EC;
defparam promx9_inst_30.INIT_RAM_1B = 288'hCAE572B95CAE572B95CAE572B95CAE572B95BADD6EB75BADD6EB75AAD56A9549A4D226F3;
defparam promx9_inst_30.INIT_RAM_1C = 288'hBADD6EB75BADD6EB75AAD56A95489A89A6F39A552A975BADD6EB75BAE572B95CAE572B95;
defparam promx9_inst_30.INIT_RAM_1D = 288'hBADD6EB75BAE572B95CAE572B95CAE572B95CAE572B95CAE572B75BADD72B5489C216554;
defparam promx9_inst_30.INIT_RAM_1E = 288'h32A150A864309A4764B248F4886532154CA6533198F075300F48A25132B5C506944E6954;
defparam promx9_inst_30.INIT_RAM_1F = 288'hCAEDB6DB6DB6DB6DB6DB6DB6DB6DB6572B95BA8390F2A2793CDE2D33E101A8642A190C86;
defparam promx9_inst_30.INIT_RAM_20 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6D95BAAC4512592D1A4B2592C968D26B30C2EBB5CAE572B95;
defparam promx9_inst_30.INIT_RAM_21 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_22 = 288'h50A05C50261B42A975CAE572B95CAE572B95CAE576BB6DAE5B2B96DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_23 = 288'h8A451E6F3691C9CC85C098A4763D250F49A3D260F0784508870942A1E12050281409C2A1;
defparam promx9_inst_30.INIT_RAM_24 = 288'hCAE572B95CAE572B95CAE572B95BADD72B95CAE572B95BADD6EB75BADD6EB75AAD52A934;
defparam promx9_inst_30.INIT_RAM_25 = 288'h58B222754BADD6EB75BADD6EB75AAD56A93489A89E6F39A4D2A954BADD6EB75BADD6EB95;
defparam promx9_inst_30.INIT_RAM_26 = 288'h79CD2A955BADD6EB75BAE572B95CAE572B95CAE572B95CAE572B95BAE56EB75BADD6EB54;
defparam promx9_inst_30.INIT_RAM_27 = 288'h42A154C8553214CA86432160E85432150A86433194CC663B1A0E03F1D1144E364EB460B2;
defparam promx9_inst_30.INIT_RAM_28 = 288'hCAE572B95DB6DB2DB6DB6DB6DB6DB6572BB6CAE572AF243A1F584F27EAD0AA6C1A9FDA86;
defparam promx9_inst_30.INIT_RAM_29 = 288'hDB6DB6DB6DB6DB6BB6DB6DB6DB6DB6DB6DB6CAE56A89165E9F9166A349ACC498A5D72BB6;
defparam promx9_inst_30.INIT_RAM_2A = 288'hCB65B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_2B = 288'h9140A050260A854320D2B8D8B52CB6532B75CAE572B95CAE572B95DAED72DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_2C = 288'hAA552691489BCDA6D238F3A0D2131D12C7648169309A4D26134983B2B87C2C1A158EC7E5;
defparam promx9_inst_30.INIT_RAM_2D = 288'hBADD72B95CAE572B95CAE572B95CAE572B95CADD72B95CAE56EB75BADD6EB75BADD6AB55;
defparam promx9_inst_30.INIT_RAM_2E = 288'hBADD6EB348542A2975BADD6EB75BADD6EB75AAD52693489A8DE7139A552A975BADD6EB75;
defparam promx9_inst_30.INIT_RAM_2F = 288'hD694164F39A4D2AB75BADD6EB95CAE572B95CAE572B95CAE56EB75CAE572B95CADD6EB75;
defparam promx9_inst_30.INIT_RAM_30 = 288'h91796528532A154CA6532954CA64331D4EA6532194CA6532994CC663B9C07A36120ACAAA;
defparam promx9_inst_30.INIT_RAM_31 = 288'hCAE576BB6CAE572B95CAEDB2B95CAEDB6DB6CAE572B95CADD48E87437309E2F63A14CBE4;
defparam promx9_inst_30.INIT_RAM_32 = 288'hDB6DB6DB6DB6DB6DB5DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D72B95BACD226D26944E6995;
defparam promx9_inst_30.INIT_RAM_33 = 288'hCB6DB6DB6CB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_34 = 288'h00C92C763A179605228138942C4A08030B2382D52E995CAE572B95CAE572B95CAED72BB6;
defparam promx9_inst_30.INIT_RAM_35 = 288'hBAD56AB54AA4D2691379B4D647107C19408491C8EC6E2C269309A4C1E92C7A450B8943A2;
defparam promx9_inst_30.INIT_RAM_36 = 288'hBADD6EB75BADD72B95CADD72B95CAE572B95CAE572B75CAE572B75CAE56EB75BADD6EB75;
defparam promx9_inst_30.INIT_RAM_37 = 288'hCAE56EB75BADD6AB3463FBAA975BADD6EB75BADD6AB55AA552A93469289A7139A552A975;
defparam promx9_inst_30.INIT_RAM_38 = 288'h4101DD78D182C9E7149A4D2AB75BADD6EB75CAE572B95CAE572B95CAE572B95BAE56EB75;
defparam promx9_inst_30.INIT_RAM_39 = 288'h4311984E371C8CCC86432190CA6532994CE753299CEA6432990CA6533194CC66381388A2;
defparam promx9_inst_30.INIT_RAM_3A = 288'hCAE576D95DAED72BB6BAE572B95CAE5B2B95CAE572BB6CAE572B958991C8A4543DADD286;
defparam promx9_inst_30.INIT_RAM_3B = 288'hDAED76DB6DB6DB6DB6DB6DB6DB6DB6D76DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6572B95;
defparam promx9_inst_30.INIT_RAM_3C = 288'hCAE576BB6DB6572DB6DB6DB6DB6DB6DB6DB6DB6DB6DD6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_30.INIT_RAM_3D = 288'h61B0D86A340E080184B1E0E85E581409C4A1405078441C2C8FD594CADD6EB95CAE572B95;
defparam promx9_inst_30.INIT_RAM_3E = 288'hBADD6EB55AAD56A9349A4D226F369AC92231A3D8508A181592C783D269309A4C260F08A0;
defparam promx9_inst_30.INIT_RAM_3F = 288'h9A4D2A975BADD6EB75BADD6EB75CAE56EB95CAE572B75CAE572B95CADD72B75BADD6EB75;

pROMX9 promx9_inst_31 (
    .DO({promx9_inst_31_dout_w[26:0],promx9_inst_31_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_37),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_31.READ_MODE = 1'b1;
defparam promx9_inst_31.BIT_WIDTH = 9;
defparam promx9_inst_31.RESET_MODE = "SYNC";
defparam promx9_inst_31.INIT_RAM_00 = 288'hCADD72B75BAE56EB75BADD6E8F274A46A955BADD6EB75BADD6EB55AA552693407B8DA713;
defparam promx9_inst_31.INIT_RAM_01 = 288'h4379504A22442F1A30593CE2934AA556EB75BADD6EB75BAE572B95CAE572B95CAE56EB95;
defparam promx9_inst_31.INIT_RAM_02 = 288'h43BA48A458141206E472410CC65432194C8653299CEA6536910AA64321D4AA65329D4EA7;
defparam promx9_inst_31.INIT_RAM_03 = 288'hDAEDB6BB5DB6576DB6DB6572BB5CAE572B95CAE572B95CAE572B95CAE56E830339148A45;
defparam promx9_inst_31.INIT_RAM_04 = 288'hDB6DB6DB6DB6DB6DB6DB6DB6BB6DB6D76DB6DB6DB6DB6DB6D76BB6DB6DB6DB6DB6DB6DB5;
defparam promx9_inst_31.INIT_RAM_05 = 288'hCAE572B95CAE572B95CAE572D96CB65B6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_31.INIT_RAM_06 = 288'hD1D8EC2A36130D86A220A8D03C210F1707638171244E2F12894480F1987090457E532B95;
defparam promx9_inst_31.INIT_RAM_07 = 288'hBADD6EB75BADD6EB55AAD5269348A44DE6D359248A2C631F8D0323B269749A4E26930983;
defparam promx9_inst_31.INIT_RAM_08 = 288'h043B1A7139A4D2A955BADD6EB75BADD6EB75BAE572B75BAE572B75BADD6EB75BADD6EB75;
defparam promx9_inst_31.INIT_RAM_09 = 288'hCAE572B75BADD6EB75BADD6EB75BAD56A84F852CAA955BADD6EB75BADD6AB54AA5526913;
defparam promx9_inst_31.INIT_RAM_0A = 288'h5331D4C8612A05044985E3460B169C526934AA556EB75BADD6EB75CADD72B95CAE572B95;
defparam promx9_inst_31.INIT_RAM_0B = 288'h229148A45640984A067238DC84881E14CC4542A190C86532990D08712990C86431994CA7;
defparam promx9_inst_31.INIT_RAM_0C = 288'hDB6DB6DB6DB6DB6BB6DB6DB6DB6DB6D76B95CADD72B95CAE572BB6CAE572B95CADD01E66;
defparam promx9_inst_31.INIT_RAM_0D = 288'hDB6DB6DB6DAEDB6DB6DB6D76DB6DB6DB6DB5DAED76DB6DB6DB6DB6DB6DB6DB6DB6DB6DB5;
defparam promx9_inst_31.INIT_RAM_0E = 288'hB249AE775CAE572B95CAE572B95CAE572BB6CB65B6BB5DB6DB2DB6DB6DB6DB6DB6DB6DB6;
defparam promx9_inst_31.INIT_RAM_0F = 288'hE26938984C210D44C251B09864151A8D44C34070883A5B1D8E03A481A0944C251D8BC421;
defparam promx9_inst_31.INIT_RAM_10 = 288'hCADD6EB75BADD6EB75BADD6EB55AA55269348A3CDE6D2491C40D2471186C984D250F49C4;
defparam promx9_inst_31.INIT_RAM_11 = 288'hAA4D2691381AC9A7139A552A954BADD6EB75BADD6EB75CADD6EB75CADD72B95CADD6EB75;
defparam promx9_inst_31.INIT_RAM_12 = 288'hBAE572B95BAE572B75BADD6EB75BADD6EB75BAD52692AA5B4AA955AADD6EB55BAD56A954;
defparam promx9_inst_31.INIT_RAM_13 = 288'h32A190DE5532194C8612A074CEBC6FBCE2D289CD26954AA556EB75BADD6EB75CAE56EB75;
defparam promx9_inst_31.INIT_RAM_14 = 288'hBA8C04A46229188C2512895C4E371B8DC8E361C12CA05329950CA6532998EA7914118C65;
defparam promx9_inst_31.INIT_RAM_15 = 288'hDB6DB6DB6DAEDB6DB6DB6D76BB5DB6D76BB5DAE576BB5BADD72B95CAE572B95BAE56EB74;
defparam promx9_inst_31.INIT_RAM_16 = 288'hDB6DB6DB6DB6D76DB5DB6DB6DB6DAEDB6BB6DB6D76DB6DB6D76DB6DAEDB6DB6DAEDB6DB6;
defparam promx9_inst_31.INIT_RAM_17 = 288'h31206C963C110DC925BADD2EB95CAE572B95CAE572B95CAED76BB5DAEDB6BB5DB6DB6DB6;
defparam promx9_inst_31.INIT_RAM_18 = 288'h70E9389C4E269347A4C2A8586C361A8882A261A8944A34120901A251E9349848148F4481;
defparam promx9_inst_31.INIT_RAM_19 = 288'hCAE56EB75BADD6EB75BADD6EB75BAD56AB54AA4D2691489BCDA4923883E4B6132289C543;
defparam promx9_inst_31.INIT_RAM_1A = 288'hBAD52A954AA4D26913512C9E7139A552A954BADD6EB75BADD6EB75BADD6EB75BAE56EB75;
defparam promx9_inst_31.INIT_RAM_1B = 288'hBADD6EB75CAE56EB75BAE56EB95BADD6EB75BADD6EB75AA5522687F7BCE6954BAD56EB75;
defparam promx9_inst_31.INIT_RAM_1C = 288'h23C120903E221CCD64532990C6612A840F0BD70C162F38A4D26954AAD52EB75BADD6EB75;
defparam promx9_inst_31.INIT_RAM_1D = 288'hBADD6EB7579E108A25229148A45E2B8E08E28238DC6E371B8E06C3E2918CC86639950CA7;
defparam promx9_inst_31.INIT_RAM_1E = 288'hDAED76DB5DAED76DB6DB6DB6DB6DB6D76DB6CAEDB6BB6CAED72BB5CAE572B95CAE572B95;
defparam promx9_inst_31.INIT_RAM_1F = 288'hDB6DB6DB6DB6DB6BB6DB6DB6DB5DAED72BB5DB6D76DB5DAEDB6BB5DAED76BB5DB6D76B95;
defparam promx9_inst_31.INIT_RAM_20 = 288'hC1C0E84E2B0A068964C281EC8C2927AEE954CAE572B95CAE572B95CAED72B95DAED76BB5;
defparam promx9_inst_31.INIT_RAM_21 = 288'h41D130943E271389C5E269349A55030D86C361A08C2C35128986A220B0946A23070A0983;
defparam promx9_inst_31.INIT_RAM_22 = 288'hBADD6EB75BADD6EB75BADD6EB75BADD6EB75AAD56A9549A4D2271379B49647128F11CDC3;
defparam promx9_inst_31.INIT_RAM_23 = 288'hAA556EB55AAD52A954AA4D268D261AC9E7349A552A975BADD6EB75BADD6EB75BADD6EB75;
defparam promx9_inst_31.INIT_RAM_24 = 288'hBADD6EB75BADD6EB95CADD72B95CADD6EB75BADD6EB75BADD6EB75AA55226C8183CE6954;
defparam promx9_inst_31.INIT_RAM_25 = 288'h331994F048238E070482412070412A9D0C8612A880F4CE7141A4F38A4D2A954BADD6EB75;
defparam promx9_inst_31.INIT_RAM_26 = 288'hCAE572B75BADD6EB34E338F0845229144CE38238F4A4771B8D86C371B8DC72475C0F0887;
defparam promx9_inst_31.INIT_RAM_27 = 288'hDAEDB2BB6CAED76D95DB6D76BB5DB6DB6DB6DB6DB6BB6DB6DB6BB5CAE572B95CAE56EB95;
defparam promx9_inst_31.INIT_RAM_28 = 288'hCAE572B95DB6D76BB5DB6DB6BB5CAED76BB5DAED72BB5DAED76DB5DAED76BB5CAED76BB5;
defparam promx9_inst_31.INIT_RAM_29 = 288'h512090161A26130763B1C8FC4A1A261B4B656129208F0BAE572B95CAE572B95CAE572B95;
defparam promx9_inst_31.INIT_RAM_2A = 288'hE749EC66230B8DC563F2F178BC4E2F17496161B0D86C36190586A251289444161A8986A2;
defparam promx9_inst_31.INIT_RAM_2B = 288'hBADD6EB75BADD6EB75BADD6EB75BADD6EB75BAD56AB55AAD52A9349A4D228F369AC92271;
defparam promx9_inst_31.INIT_RAM_2C = 288'h283CE6934AA552A954AA552A954AA4D2268AC334A27139A552A954BADD6EB75BADD6EB75;
defparam promx9_inst_31.INIT_RAM_2D = 288'hAA552EB75BADD6EB75BADD6EB95CADD6EB75BADD6EB75BADD6EB75BADD6EB55AA4D1A709;
defparam promx9_inst_31.INIT_RAM_2E = 288'h71C930AEA926944CC28238E0904824120703332994C86022880F4CF79C5A4F39A4D2A955;
defparam promx9_inst_31.INIT_RAM_2F = 288'hBAE572B75CAE572B75BADD6E89161B8DC74322899C6E48191C8A4681B124B259230E08E3;
defparam promx9_inst_31.INIT_RAM_30 = 288'hCAE576B95CAED72B95CAE572B95DAED76BB5CAED76B95DB6572B95CAE572B95CAE576D95;
defparam promx9_inst_31.INIT_RAM_31 = 288'hCAE572B95CAE572B95CAED76BB5DAED72BB5DAED76BB5CAED76BB5CAED76B95DAE572B95;
defparam promx9_inst_31.INIT_RAM_32 = 288'h61B0D44A230A0586A240806C983C1D8F070332B0A06E3D3409074372DCF2D95CAE572B95;
defparam promx9_inst_31.INIT_RAM_33 = 288'h69248E230E21918662F1D9309848150F8BC5F281608A261B0D86A220B0D86C361A88C2A2;
defparam promx9_inst_31.INIT_RAM_34 = 288'hBADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6AB55AAD5269349A45226F3;
defparam promx9_inst_31.INIT_RAM_35 = 288'hAA4D1A4E938C4E6934AA552A954AA552A9549A4D226C328B4A27349A552A954BADD6A954;
defparam promx9_inst_31.INIT_RAM_36 = 288'h9A4D2A955BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6AB54;
defparam promx9_inst_31.INIT_RAM_37 = 288'h82C968AE39240DC765920A2890382412090471B91C72443A9D0C6512B0B8D6CF7A45A513;
defparam promx9_inst_31.INIT_RAM_38 = 288'hCAE572B95BADD6EB75BAE56EB75BAD5268495130D86E481B8DC7E623114CC46924964B25;
defparam promx9_inst_31.INIT_RAM_39 = 288'hDAE576B95DAE572BB5CAE572B95DAE572B95DAE572BB5DAE576B95DB6572BB5DAE572B95;
defparam promx9_inst_31.INIT_RAM_3A = 288'hBAE532B95CAE572B95CAE572B95CAE576B95DAE576B95CAE572B95CAE576BB6DAE576B95;
defparam promx9_inst_31.INIT_RAM_3B = 288'h61A8904C361B0D86C330B0D84C25138EC963B1E930763A130F82E2E39A7D14392C8E4F74;
defparam promx9_inst_31.INIT_RAM_3C = 288'h9A45226F369244A1CE8250D4482917178BA4D26920523F2E9544C25128944825130D86C3;
defparam promx9_inst_31.INIT_RAM_3D = 288'hBAD52A975BADD6EB75BADD72B75BADD6EB75BADD6EB75BADD6EB55AADD6AB55AACD26934;
defparam promx9_inst_31.INIT_RAM_3E = 288'hAAD56AB54AA44F9B2A48C4E2934AA552A954AA55269349A4D1E6C2593CE2714AA552A954;
defparam promx9_inst_31.INIT_RAM_3F = 288'hF7A45A5139A552A975AA5D6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB55;

pROMX9 promx9_inst_32 (
    .DO({promx9_inst_32_dout_w[26:0],promx9_inst_32_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_39),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_32.READ_MODE = 1'b1;
defparam promx9_inst_32.BIT_WIDTH = 9;
defparam promx9_inst_32.RESET_MODE = "SYNC";
defparam promx9_inst_32.INIT_RAM_00 = 288'h92D164B0592C964B24A2D15C6E3C2B8DC90382412090482412092413A190C66022078D6C;
defparam promx9_inst_32.INIT_RAM_01 = 288'hCAED72B95CAE572B95BADD6EB75BADD6EB75AA55227A671B0D86E371B908E25231188FE5;
defparam promx9_inst_32.INIT_RAM_02 = 288'hCAE572B95DAE572B95DAE572BB5CAE572B95DAED76BB5DB6572BB5DAE576BB5CAE572BB5;
defparam promx9_inst_32.INIT_RAM_03 = 288'hB2B834D03065D72B95CAE572B95CADD72B95CAE572B95DAE572B95DAE572B95CAE576BB6;
defparam promx9_inst_32.INIT_RAM_04 = 288'h61B0D86A26190586C361A89444161B0986A3A0E0F4783B1D8F4984B1D930724A11A51289;
defparam promx9_inst_32.INIT_RAM_05 = 288'h9A4D269348A44DE6D3591C420C172B8905C2C27178BC5E2F178B8491E0102A351A8D4461;
defparam promx9_inst_32.INIT_RAM_06 = 288'h9A552A954AA552A975BADD6EB75BADD6EB75BADD6EB75BADD6EB75BAD56EB55AAD56AB54;
defparam promx9_inst_32.INIT_RAM_07 = 288'hBADD6EB75BAD52A954AA44D518C48BCE29349A4D2A954AA4D269349A44CA0C3593CE2734;
defparam promx9_inst_32.INIT_RAM_08 = 288'h02A040F6D07A45E5139A552A954AA552EB75BADD6EB75BADD6EB75BADD6EB75BADD6EB75;
defparam promx9_inst_32.INIT_RAM_09 = 288'h239180B4592C964B2592C964B2592D940DA5A238E06E38241208E3824120904D29950E45;
defparam promx9_inst_32.INIT_RAM_0A = 288'hCAE572B95CAE572B95CAE572B95BADD6EB75BADD6EB75AA5D1A50361B0D86E371C120723;
defparam promx9_inst_32.INIT_RAM_0B = 288'hCAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAED72B95CAE572B95CAE576B95;
defparam promx9_inst_32.INIT_RAM_0C = 288'hA1512C449449A686C1B2B922575CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95;
defparam promx9_inst_32.INIT_RAM_0D = 288'h4030C82C361B0D86C320B0D86C361B0CC2A261B098640D2F8F49A4C1D8F09A4D268F0963;
defparam promx9_inst_32.INIT_RAM_0E = 288'hBAD56A955AA4D2691489BCDE6D259147DE44D1A08C323E36978BC5E2F178BC5D2E130843;
defparam promx9_inst_32.INIT_RAM_0F = 288'h5944E27349A552A954AA552A975BADD6EB75BADD6EB75BADD6EB75BADD6EB75BADD6AB75;
defparam promx9_inst_32.INIT_RAM_10 = 288'hBADD6EB75BADD6EB55AAD52A9549A44D0E716944E29349A4D2A954AA4D269349A3CDC70C;
defparam promx9_inst_32.INIT_RAM_11 = 288'h921990C4602A89138D08245E7149A552A954AA5D6EB75BADD6EB75BADD6EB75BADD6EB75;
defparam promx9_inst_32.INIT_RAM_12 = 288'h71B9209048240E0966A35164B24A2D9A8B25A2D148C46231948EE38238DC704823920904;
defparam promx9_inst_32.INIT_RAM_13 = 288'hCAE572B95CAE572B95CAE572B95CAE572B95BADD6EB75BADD6EB54AA4D162C271B8DC6E3;
defparam promx9_inst_32.INIT_RAM_14 = 288'hCAE572B95CAE56EB95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95;
defparam promx9_inst_32.INIT_RAM_15 = 288'hD269349C4C258E8764D20A1520771486C948BADD6EB74BADD6EB75CAE572B95CAE572B95;
defparam promx9_inst_32.INIT_RAM_16 = 288'h713878BC4E2B0880C26228D86A24130D86C361B0CC2C361B0CC565E271389A4E260F49A4;
defparam promx9_inst_32.INIT_RAM_17 = 288'hBADD6AB55AAD52A954AA4D2691489BCDA6B2489439CC5A1A0CCB64E3717CDE6F37978DC5;
defparam promx9_inst_32.INIT_RAM_18 = 288'h89BCD44716944E2734AA552A954AA552A975BADD6EB75BADD6EB75BADD6EB75BADD6EB74;
defparam promx9_inst_32.INIT_RAM_19 = 288'hBADD6EB75BAD56EB55BADD6A955AAD52A9549A3CD90B26944E69149A4D269349A4D26934;
defparam promx9_inst_32.INIT_RAM_1A = 288'h824120904924908E25E2A8995AE182C9E7139A552A954BADD6EB75BADD6EB75BADD6EB75;
defparam promx9_inst_32.INIT_RAM_1B = 288'h7238DC6E371C11C70482411C9038240E090481C0DC6E48239288A8439980D04824120904;
defparam promx9_inst_32.INIT_RAM_1C = 288'hCAE572B95CAE572B95CAE572B95CAE572B95CAE572B95BADD6EB75BADD6EB54AA4D1A4E3;
defparam promx9_inst_32.INIT_RAM_1D = 288'hCAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95;
defparam promx9_inst_32.INIT_RAM_1E = 288'hB1F1389C4E271389A4D26930984C1E1788273450D87818272AA975BAF3A9975BADD6EB75;
defparam promx9_inst_32.INIT_RAM_1F = 288'hF379BCD43E2F174B22F2E97C943A028D864161B0D86C36188186C361B0EC3C3F279389A4;
defparam promx9_inst_32.INIT_RAM_20 = 288'hBADD6EB74AA556AB54AA552A9549A4D2691489BCDA6B2488C35D0852215C6E2D2F178BE6;
defparam promx9_inst_32.INIT_RAM_21 = 288'h9A4D2693489AC54491693CE69349A552A954AA552A975BADD6EB75BADD6EB75BADD6EB75;
defparam promx9_inst_32.INIT_RAM_22 = 288'hBADD6EB75BADD6EB55BADD6EB55AAD56AB54AA55269349A3CDD2916944E69349A4D26934;
defparam promx9_inst_32.INIT_RAM_23 = 288'h824120904824120924824968826A2289D7AE182C9E7139A552A954BADD6EB75BAD52EB75;
defparam promx9_inst_32.INIT_RAM_24 = 288'hAA551A4078238DC6E371C1209048241208E482411C90472412090482412092491A220703;
defparam promx9_inst_32.INIT_RAM_25 = 288'hCAE572B95CAE572B95CAE572B95CAE572B95CAE572B95BADD72B95BADD6EB75BADD6EB54;
defparam promx9_inst_32.INIT_RAM_26 = 288'hBADD6EB75BAE572B95CAE572B95CAE572B95CADD6EB95CADD72B95CAE572B95CAE572B95;
defparam promx9_inst_32.INIT_RAM_27 = 288'hF2F1389A4F2F93CBE4F2713C9C4E271389C4C1E92478452E9090A250991CC8F89A89C775;
defparam promx9_inst_32.INIT_RAM_28 = 288'h61697CC06F3716C722F2F1AC9E5E2C8BCBC5E2E13426061B0944A230B0DC4C3619038BE5;
defparam promx9_inst_32.INIT_RAM_29 = 288'hBADD6EB75BADD6EB75BAD52AB55AAD52A9549A4D2693489BCDA6B2388C35D2A6318C84A3;
defparam promx9_inst_32.INIT_RAM_2A = 288'h9A4D269349A4D2691389F1C0E9169BCE69349A552A954AA552A975BAD52EB75BADD6EB75;
defparam promx9_inst_32.INIT_RAM_2B = 288'hBAD52EB75AAD56AB54AA556EB75AAD56AB55AAD52AB54AA5526934898B9927179C4E6934;
defparam promx9_inst_32.INIT_RAM_2C = 288'h8241209048241209048241209249249249025138E19CE2834A2734AA552A954AA5D6A975;
defparam promx9_inst_32.INIT_RAM_2D = 288'hBADD6EB54AA4D2264871B8DC6E382411C70471C120904824120904824120904824120904;
defparam promx9_inst_32.INIT_RAM_2E = 288'hCAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CADD72B95BADD6EB75;
defparam promx9_inst_32.INIT_RAM_2F = 288'h50B0A4975BADD6EB75BADD6EB75BADD6EB95CAE572B95CAE572B95BAE56EB95CAE572B95;
defparam promx9_inst_32.INIT_RAM_30 = 288'h41597C805F2F97C983F2F97CBE5F2F97CBE4F2713C9C4E26930984A120E88A55038C0184;
defparam promx9_inst_32.INIT_RAM_31 = 288'h74294C66161A8A89E5E2D0E4584A150E87850379BCB22F2F940BA41090146A24130D86C2;
defparam promx9_inst_32.INIT_RAM_32 = 288'hBADD6EB75BADD6EB75BADD6A955BAD52AB55AA552A9349A4D2691489BCDE6B2388C35D4C;
defparam promx9_inst_32.INIT_RAM_33 = 288'h79C4E69349A4D269349A4D229136928CA0B279C4E69349A4D26954AA552A955AA5D6EB75;
defparam promx9_inst_32.INIT_RAM_34 = 288'hAA5D6A954BADD6EB55AADD6A975BAD56AB55AAD56A954AAD52A954AA552693499A1F5AB1;
defparam promx9_inst_32.INIT_RAM_35 = 288'h824120904824120904824120904824124925A2491C704510A2DBEF48BCE2734AA552A954;
defparam promx9_inst_32.INIT_RAM_36 = 288'hBADD6EB75BADD6EB54AA4D226709238D86E3824120904824120904824120904824120904;
defparam promx9_inst_32.INIT_RAM_37 = 288'hBAE572B95CAE572B95CAE572B95CADD72B95CAE572B95CADD72B95CADD72B95CAE56EB75;
defparam promx9_inst_32.INIT_RAM_38 = 288'h735A2122051286C911AA5D6A974BADD6EB75BADD6EB75CAE56EB95CAE572B95CADD72B95;
defparam promx9_inst_32.INIT_RAM_39 = 288'h51B0D84A3A08140A05F2816C7E502817CA25F2817CBE5F2F97C9E4F26934983B1A050301;
defparam promx9_inst_32.INIT_RAM_3A = 288'h488439D4C85A9948624118606E2A1D0AC6E280C060302A150B8A05F350F4806037910460;
defparam promx9_inst_32.INIT_RAM_3B = 288'hBAD52EB54BAD52EB75AA5D6EB75BAD52A954AA552A954AA552A9349A4D269348A44DA4B2;
defparam promx9_inst_32.INIT_RAM_3C = 288'h89B2162B179C4E69149A4D269349A44E271348A88E2D279C5269349A552A954BA552A975;
defparam promx9_inst_32.INIT_RAM_3D = 288'hAA552A954AA5D6A954AA552EB54AA556A954AA556EB55BAD52A954AAD52A954AA4D26934;
defparam promx9_inst_32.INIT_RAM_3E = 288'h92412090482412090482492492482412092492412CBC79249186C35132B5C105944E6934;
defparam promx9_inst_32.INIT_RAM_3F = 288'hBAE56EB95BADD6EB75BADD6EB54AA55268F354A0586E381C120904824120924824120904;

pROMX9 promx9_inst_33 (
    .DO({promx9_inst_33_dout_w[26:0],promx9_inst_33_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_41),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_33.READ_MODE = 1'b1;
defparam promx9_inst_33.BIT_WIDTH = 9;
defparam promx9_inst_33.RESET_MODE = "SYNC";
defparam promx9_inst_33.INIT_RAM_00 = 288'hCAE56EB75CAE56EB95CAE572B95CAE572B95CAE572B95BADD72B75CAE572B95CAE572B95;
defparam promx9_inst_33.INIT_RAM_01 = 288'hC2208C48231206C3246160902A182CA6A775AADD6EB75BADD6EB75CADD72B75CADD72B75;
defparam promx9_inst_33.INIT_RAM_02 = 288'hD2F17CBE4614054480020140A05F2F100A26130140A05028140A05F2F1389E5F27134984;
defparam promx9_inst_33.INIT_RAM_03 = 288'h8A44DE6D2489439D6D963A54C84311894503A240BCAC181386030180C0A4542A1713CB64;
defparam promx9_inst_33.INIT_RAM_04 = 288'hAA552A975AA552A975BADD6A975AA5D6EB75AA5D6EB54AA552A9549A552A9349A4D26934;
defparam promx9_inst_33.INIT_RAM_05 = 288'h9A4D269337942962D279C4E27139A4D2693489C4E26F3920A162F389C5269349A5526954;
defparam promx9_inst_33.INIT_RAM_06 = 288'h79C4E6934AA552A954BAD52EB54AAD52A954AA552A954AA552A954AA552A954AA552A934;
defparam promx9_inst_33.INIT_RAM_07 = 288'h82492490492412090482412492482412090482412492492D174DAEB29868AA214533DE71;
defparam promx9_inst_33.INIT_RAM_08 = 288'hBAE56EB75BADD6EB75BADD6EB75BADD6EB54AA5526913590A144C371B8E0904824120924;
defparam promx9_inst_33.INIT_RAM_09 = 288'hBAE56EB95BADD6EB95BADD72B75CADD72B95BAE572B75CAE56EB95CAE56EB75CAE56EB95;
defparam promx9_inst_33.INIT_RAM_0A = 288'hF2F1389A431A8D84C230988C2A23058608A221B0944A499552EB75AADD6EB75BADD6EB75;
defparam promx9_inst_33.INIT_RAM_0B = 288'h8148A8583F2D8EC605F2F96C923028144A05137104A26128984C06028140A0502F97CBE5;
defparam promx9_inst_33.INIT_RAM_0C = 288'h9A4D269348A44DE6D2491C461CEB642D526732988C48230C93098371591C50180C060501;
defparam promx9_inst_33.INIT_RAM_0D = 288'h9A4D26954AA552A954BAD52A974AA5D6A954AA552EB54AA552A954AA552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_0E = 288'hAA552A9349A4D26934D63A962F269C4E27349A4D269348A44DE6F3510C162F289C526934;
defparam promx9_inst_33.INIT_RAM_0F = 288'h656B4A0D289C4E6954AA552A954AA5D6E954AA552A954AA552A954AAD56A954AA552A954;
defparam promx9_inst_33.INIT_RAM_10 = 288'h92412492492492492482492490492412492482492490492492494504536CA0820A0904E3;
defparam promx9_inst_33.INIT_RAM_11 = 288'hBADD72B95CAE572B75BADD72B75BADD6EB75AAD56EB54AA4D2691379AC490815130DC704;
defparam promx9_inst_33.INIT_RAM_12 = 288'hBADD6EB75BADD72B95BAE572B95CAE56EB75BAE572B95CADD72B95CAE572B95CAE56EB75;
defparam promx9_inst_33.INIT_RAM_13 = 288'h02817CBE5F2713898391A89C68251289448130A08C281B0B10836461A92A975BADD2E975;
defparam promx9_inst_33.INIT_RAM_14 = 288'hE3616470280C060322A150B096471613CBE5B1D8FCA05B18144C26130984C25028144C05;
defparam promx9_inst_33.INIT_RAM_15 = 288'hAA552A9549A4D2693489C4DE6F369248A20FD74B2168A41180468382985C784A1E9607A6;
defparam promx9_inst_33.INIT_RAM_16 = 288'h89CD269349A4D2A9549A552A954AA552A954AA552E954AA552A954AA552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_17 = 288'hAA552A954AA55269349A4D228F333FB922D279C4E27149A4D2691489C4DE6305114164F3;
defparam promx9_inst_33.INIT_RAM_18 = 288'h30A8904AAC68C164D289CD26954AA552A954BA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_19 = 288'hD320944C372412CACA03D16492492492492492412492482412492492C968A8AB6DB58661;
defparam promx9_inst_33.INIT_RAM_1A = 288'hBADD6EB75BADD6EB75BADD72B75BADD6EB75BADD6EB75BADD6EB54AA552693489BCD63EF;
defparam promx9_inst_33.INIT_RAM_1B = 288'hAA556EB74BA5D6EB75BADD6EB75BADD6EB95CADD72B75CADD6EB75CAE56EB75CADD72B75;
defparam promx9_inst_33.INIT_RAM_1C = 288'h130984C2512817CBE5F2F13876651C930AC3824920924612890463412854B64B1C0D43AA;
defparam promx9_inst_33.INIT_RAM_1D = 288'h9259688C271F1F4DA7E338A43025130401048171685C503796C702028984C46130944C26;
defparam promx9_inst_33.INIT_RAM_1E = 288'hAA552A954AA552A9549A4D269349A44E26F3692492230F7EBA58CB761874C4032B92CCC3;
defparam promx9_inst_33.INIT_RAM_1F = 288'h75A4564F389CD269349A4D2A954AA552A954AA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_20 = 288'hAA552A954AA55269349A4D269349A4D228D26424522D279C4E27148A452271489C4DA4A2;
defparam promx9_inst_33.INIT_RAM_21 = 288'h51184C24051289554C07A45E6F389CD26954AA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_22 = 288'h89BCDE6B138A2646A251B0E498D34B2C93CE03E3A8B2492492092492492492465DB78FAE;
defparam promx9_inst_33.INIT_RAM_23 = 288'hBADD6EB75BADD72B75BADD6EB75BADD6EB95BADD6E975BADD6EB75AAD56EB75AA5526934;
defparam promx9_inst_33.INIT_RAM_24 = 288'hB250E468121D4EA955AA5D6EB75BADD6EB75BADD72B75BADD6EB75BADD72B75BADD6EB95;
defparam promx9_inst_33.INIT_RAM_25 = 288'h130984C26130984C2602817CBE5F2F13494361E1B0D86A2C92CB6592516490340A084143;
defparam promx9_inst_33.INIT_RAM_26 = 288'h519810988C41858523C2B89C72462580404130984C2821039645E5817100C26130984C25;
defparam promx9_inst_33.INIT_RAM_27 = 288'hAA552A954AA552A954AA552A9349A4D269349A4D226F369AC96471187BF1D2C652290565;
defparam promx9_inst_33.INIT_RAM_28 = 288'h79BCD648207AC9A4F389CD229349A4D26934AA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_29 = 288'hAA552A9549A552A954AA55269349A4D269348A44DE7A6B21C522B279BCE271389C522713;
defparam promx9_inst_33.INIT_RAM_2A = 288'hD3698C4613098586A251226D9EF48B49E7139A4D26954AA552A954AA552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_2B = 288'hAA552A9349A44E26F3592445E079228944C3820A196AAE78A28B6D75CB11565B2EBA9B4D;
defparam promx9_inst_33.INIT_RAM_2C = 288'hBADD72B75BADD6EB75BADD6EB75BADD2EB75BADD6EB74BADD6E975BAD56A975BADD6EB54;
defparam promx9_inst_33.INIT_RAM_2D = 288'hA238C4146B1D928943509095F74AA5D6E975BADD6EB75BADD6EB75BADD32B75BADD6EB75;
defparam promx9_inst_33.INIT_RAM_2E = 288'h0311C4C26130984C26128984C26028140BE5F26930CC3A2E1B0D86D371FD1E8E3F1F4D86;
defparam promx9_inst_33.INIT_RAM_2F = 288'h9632945C655104D5A24249B0E8140C8F0AE480A84C26130984C26131208C2C4A1F96C7A4;
defparam promx9_inst_33.INIT_RAM_30 = 288'hAA552A954AA552A954AA4D2A954AA55269549A4D269349A4D2271379BCD64B2388C3DFAE;
defparam promx9_inst_33.INIT_RAM_31 = 288'h89C4E271379B4D54E3282C9E71389CD269349A4D2A954AA552A9549A552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_32 = 288'hAA552A954AA552A954AA552A9349A4D269349A4D2693489B4D94A220D10A0B2693CE2713;
defparam promx9_inst_33.INIT_RAM_33 = 288'hC31270D044120A888230D1144E3656341E91693CE27349A4D2A9349A552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_34 = 288'hBAD56A954AA552A9549A4D2271379B49627007B280EA261B0DC6E4925168A284573F5D86;
defparam promx9_inst_33.INIT_RAM_35 = 288'hBADD2EB95BADD6EB75BADD6EB75BADD6EB75BADD2EB75BADD6EB75BADD6A975BAD56EB75;
defparam promx9_inst_33.INIT_RAM_36 = 288'hF471F4F86A2A8D05C2A1D128743A1B88C24FBA552A974BA5D6EB74BA5D6EB75BADD6EB74;
defparam promx9_inst_33.INIT_RAM_37 = 288'h6118E87E540697CC26130984C26230984C0502817CBE5E2692C8C2C361B0DA6E3F1FD1E8;
defparam promx9_inst_33.INIT_RAM_38 = 288'h489C4600FE7636174520F9F0BC72010D04C4E420902E2E2F87066140984C26130984C2A2;
defparam promx9_inst_33.INIT_RAM_39 = 288'hAA5526954AA4D26954AA552A954AA5526954AA4D269549A4D269349A4CE271379BCDA6B2;
defparam promx9_inst_33.INIT_RAM_3A = 288'h693CDE71389C4E26F379BC947EF48AC9E71389C5269349A4D269349A4D269349A552A934;
defparam promx9_inst_33.INIT_RAM_3B = 288'hAA552A954AA4D26954AA552A954AA4D269349A4D269349A452291379B49C661416341E91;
defparam promx9_inst_33.INIT_RAM_3C = 288'h71B924945B2D94C46182185456551308D32BD68C122D279C4E67349A552A954AA552A954;
defparam promx9_inst_33.INIT_RAM_3D = 288'hBADD6EB75AAD52A954AA552A954AA4D2691489BCDA4B2489C0A18D1401D86C26130DC6E4;
defparam promx9_inst_33.INIT_RAM_3E = 288'hBADD2EB75BADD6A974BADD6EB75BADD6EB75BADD6EB75BADD6EB74BADD6EB75BADD6EB75;
defparam promx9_inst_33.INIT_RAM_3F = 288'hE3F9FD1E8F3F1F4F86922890420A1D12474491C8DC66069552A954BA5D6E975BADD2E974;

pROMX9 promx9_inst_34 (
    .DO({promx9_inst_34_dout_w[26:0],promx9_inst_34_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_43),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_34.READ_MODE = 1'b1;
defparam promx9_inst_34.BIT_WIDTH = 9;
defparam promx9_inst_34.RESET_MODE = "SYNC";
defparam promx9_inst_34.INIT_RAM_00 = 288'h4130E48A271A8984808271603C5131188C26130144C2613797CBE5E20098745C369F4DC7;
defparam promx9_inst_34.INIT_RAM_01 = 288'h89C4DE6D2692C92250187BF5D6D554B0824155228CA6341A0F0CA240C8B0BA170A04C4A2;
defparam promx9_inst_34.INIT_RAM_02 = 288'h9A4D2A954AA4D2A954AA4D26934AA552A934AA4D2A954AA4D269349A4D269349A4CE2714;
defparam promx9_inst_34.INIT_RAM_03 = 288'h417381E91593CDE6F379BCDE6F3692A9862F48B49E71389CD269349A4D269349A4D26954;
defparam promx9_inst_34.INIT_RAM_04 = 288'hAA5526934AA552A9549A4D26934AA552A954AA4D269349A4D269348A44E26F369AC94482;
defparam promx9_inst_34.INIT_RAM_05 = 288'h1389C9008A2D970D0340984C344F3B8D86E344C2F5A0F382C9A6F389CD26934AA4D2A954;
defparam promx9_inst_34.INIT_RAM_06 = 288'hBADD6A974AADD6A954AAD52A954AA552A954AA4D269348A44E26F3692C964711783E59A5;
defparam promx9_inst_34.INIT_RAM_07 = 288'hBADD6EB75BADD6E975BADD6A974BADD6EB75BADD6EB75BADD6EB75BA5D72B75BA656EB75;
defparam promx9_inst_34.INIT_RAM_08 = 288'hC361B4FC7E3F9FCFE8F3F1F4F86619854200A2512C944A1D0E86A4314CEA954AA552E954;
defparam promx9_inst_34.INIT_RAM_09 = 288'h9268942615130D44824128840E1311820BA5708144C26130984A0502F9789C5E32098766;
defparam promx9_inst_34.INIT_RAM_0A = 288'h9A44E27348A44DE6F379B4964913894061CFC74B1144824512CCA541A1146A3A31858584;
defparam promx9_inst_34.INIT_RAM_0B = 288'h9A4D269349A552A9549A552A934AA4D2A9549A4D269349A4D269349A4D26934AA5526934;
defparam promx9_inst_34.INIT_RAM_0C = 288'h69140C46161F3860915934DE6F379BCDE6D25928B1A3058B4DE71389CD269349A4D26934;
defparam promx9_inst_34.INIT_RAM_0D = 288'h9A4D269349A4D269549A4D269349A4D269549A552A9349A4D269349A4D2693489C4DE6F3;
defparam promx9_inst_34.INIT_RAM_0E = 288'h48A44A030F7DB5D5E6B27980FC6B240DC6A2A2225D56DE70BCE291693CE27139A4D26934;
defparam promx9_inst_34.INIT_RAM_0F = 288'hBADD6E974BADD6E954BADD6AB75AA556A954AA552A954AA55269349A452291379BCDA4B2;
defparam promx9_inst_34.INIT_RAM_10 = 288'hAA552A974BADD6EB74BADD6EB74BADD2A954BADD6EB75BADD2E974CADD6EB75BADD6EB75;
defparam promx9_inst_34.INIT_RAM_11 = 288'h7128ACB66C369B8FE7F3F9FCFE7E3F1F4D45412090441C250E8943A1D1248C8E12966954;
defparam promx9_inst_34.INIT_RAM_12 = 288'h51A8E8A817169485A361289448230A85822120A08C260A1D0EC626128984C05F2F938BA3;
defparam promx9_inst_34.INIT_RAM_13 = 288'h9A4D269349A4D2693489C4E26F379B49A6B259244E25007F3ADB0B6522490664228D46A3;
defparam promx9_inst_34.INIT_RAM_14 = 288'h9A4D269349A4D269349A4D26934AA4D2A9349A4D269549A4D26934AA4D269349A4D26934;
defparam promx9_inst_34.INIT_RAM_15 = 288'h89C4DE6F35969A488275F3860915934DE6F369B49A47131208503059349E71389CD26934;
defparam promx9_inst_34.INIT_RAM_16 = 288'h9A4D269349A4D269349A4D269549A4D26934AA55269349A4D269349A4D269349A4D26713;
defparam promx9_inst_34.INIT_RAM_17 = 288'h89C4DE6F37934964B1389C0A00FF773B1D6DA6D32DB8EE77B85E5038AC9A4F379C4E2714;
defparam promx9_inst_34.INIT_RAM_18 = 288'hBADD2A974BA552EB75BA552A954AA556AB75AAD56A954AA552A954AA55269349A4D22713;
defparam promx9_inst_34.INIT_RAM_19 = 288'h9670A1134AA552A954BA552E974BA5D6E974BA5D6E954AA5D2E974BA5D6A975BADD2EB75;
defparam promx9_inst_34.INIT_RAM_1A = 288'hF2F1348C0514128B66C369F8FE7F3FA3CFC7E3E9F0AC330A890461C25128964A1D0E47A5;
defparam promx9_inst_34.INIT_RAM_1B = 288'h91314828351A8D46A37220645A510E0D44A2D2508824130A8904E220D878AC1F28180A05;
defparam promx9_inst_34.INIT_RAM_1C = 288'h9A4D269349A4D269349A4D2693489C4E271379BCDE6D3692C96491280C01FAEB6C2D5488;
defparam promx9_inst_34.INIT_RAM_1D = 288'h89CD269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_34.INIT_RAM_1E = 288'h9A4CE271389C4DE6D248A88C2A2D77B8E291593CDE6D2692C9234C30A0A160F48B49E713;
defparam promx9_inst_34.INIT_RAM_1F = 288'h89C4E29349A4D269349A4D269349A4D269349A4D269349A552A9349A4D269349A4D26934;
defparam promx9_inst_34.INIT_RAM_20 = 288'h9A4D269348A4D2291389BCDE6F2592C9629148A44E27128140E27148AC564D2693CDE713;
defparam promx9_inst_34.INIT_RAM_21 = 288'hBA5D2EB54BAD52E975BA552E974BA5D2E954AA556AB54AAD56AB54AA552A954AA552A934;
defparam promx9_inst_34.INIT_RAM_22 = 288'hA1D124784C6EB8086EAA552A954BA5D6A975AA552A954BADD6E954AA5D6E974BA5D2A974;
defparam promx9_inst_34.INIT_RAM_23 = 288'h8150F8BE5E27128283514968B66C371F8FE8F3F9F8FC7D3E1A486130A090440A250E8744;
defparam promx9_inst_34.INIT_RAM_24 = 288'hF7E3A990B5499B84822090946A351A8D44A2A1E170282D19044282512090461414108123;
defparam promx9_inst_34.INIT_RAM_25 = 288'h9A4D269349A4D269349A4D269349A4D2691489C4E271389C4DE6F379B4964B2491C4A010;
defparam promx9_inst_34.INIT_RAM_26 = 288'h49349E71389C5269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_34.INIT_RAM_27 = 288'h9A4D2693499CCE271389BCDE6D2A62890482E704122B26934DE6D2692C4A02830A0ADA30;
defparam promx9_inst_34.INIT_RAM_28 = 288'h89C4E27138A4D269349A4D269349A4D269349A4D269349A4D269349A55269349A4D26934;
defparam promx9_inst_34.INIT_RAM_29 = 288'hAA552A9549A4D269349A4D269348A44E271379BCDA6D269B49A4D2692C9A4D3793CDE713;
defparam promx9_inst_34.INIT_RAM_2A = 288'hBA552E974AA552A954BA5D2E954AA5D2A954AA552A954AAD52A955AA552A954AA552A954;
defparam promx9_inst_34.INIT_RAM_2B = 288'hA238A0544A1D124763C773F9E4789CD26954AA552A975AA552A954BA5D2A954AA552E975;
defparam promx9_inst_34.INIT_RAM_2C = 288'h309898462E0E1245C4D270946A2A2D168B65C369FCFC7F3F1F8FC7C3599866130A094761;
defparam promx9_inst_34.INIT_RAM_2D = 288'h692C8E2712803F9D8DA63A910806228842426228D46825130586E430904C4A330984C282;
defparam promx9_inst_34.INIT_RAM_2E = 288'h9A55269349A4D269349A4D269349A4D269349A4D229348A452271389C4E26F379BCDA6D2;
defparam promx9_inst_34.INIT_RAM_2F = 288'h30D175C504934DE7138A4D229349A4D269349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_34.INIT_RAM_30 = 288'h9A4D269349A4D269349A44E271389BCDE6D26198904CA0794522D26934DA6D2592452282;
defparam promx9_inst_34.INIT_RAM_31 = 288'h79C4E271389C5269349A4D269349A4D269349A4D269349A4D269549A4D269349A4D26934;
defparam promx9_inst_34.INIT_RAM_32 = 288'hAA552A954AA552A9349A4D269349A4D269349A4D2291389C4DE6F379BCDE6F379BCDE713;
defparam promx9_inst_34.INIT_RAM_33 = 288'hAA552E975BA5D2A954BA5D2A975BAD52E954AA552A954AA552A934AA552A954AA552AB54;
defparam promx9_inst_34.INIT_RAM_34 = 288'h4120882C4A1D92894360C8E4646F7FBF5F6D44CD2A954AA552A974AA552A954BA5D2A954;
defparam promx9_inst_34.INIT_RAM_35 = 288'h30984C26131204C6A1722838AE2A03110545C2D168B45C369B4DA7E3F1F8FA7C34910482;
defparam promx9_inst_34.INIT_RAM_36 = 288'h79BCDE6D369B496491489C4E00FE75B216A92390D06822090586C451A8E46E2E3F08CC60;
defparam promx9_inst_34.INIT_RAM_37 = 288'h9A4D269349A4D269349A4D269349A4D269349A4D269349A4D229348A452271389C4E2713;
defparam promx9_inst_34.INIT_RAM_38 = 288'h59244A06130D179C705934DE71389CD269349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_34.INIT_RAM_39 = 288'h9A4D269349A4D2693499CD2673399CCE271389BCDE6B238B28D20F179C564D2793CDA6D2;
defparam promx9_inst_34.INIT_RAM_3A = 288'h89C4E271389C52691389C5269349A4D269349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_34.INIT_RAM_3B = 288'hAA552AB54AA552A954AA4D2A934AA4D2A934AA4D269349A4D269348A452271389C4E2713;
defparam promx9_inst_34.INIT_RAM_3C = 288'hAA5D2E954AA552A954AA552A954BADD2A954AA552A954AA552A954AA5526954AAD52A954;
defparam promx9_inst_34.INIT_RAM_3D = 288'hB2B0D0461412880163A2592C964A1C8E04A0E383F9DAE75A426954AA552A954AA552A954;
defparam promx9_inst_34.INIT_RAM_3E = 288'h40C084DA512205046130989048230C10C1A33028D8745A2C968B45D361B0DA7E3F1F8FA6;
defparam promx9_inst_34.INIT_RAM_3F = 288'h89C52271379C4DE6F379BCDA4B25924922712803F9D6C95AA14A834128882C46239186A2;

pROMX9 promx9_inst_35 (
    .DO({promx9_inst_35_dout_w[26:0],promx9_inst_35_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_45),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_35.READ_MODE = 1'b1;
defparam promx9_inst_35.BIT_WIDTH = 9;
defparam promx9_inst_35.RESET_MODE = "SYNC";
defparam promx9_inst_35.INIT_RAM_00 = 288'h9A4D269349A4D269348A4D269349A4D269349A4D269349A4D269349A4D2693489CD22913;
defparam promx9_inst_35.INIT_RAM_01 = 288'h79BCDE4D259247DE41309A7DE91693CDE71389CD227349A4D269349A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_02 = 288'h9A4D269339A4D269349A4D2693499CD2693499CCE271389C4DE6D269244E27148AC9A4F2;
defparam promx9_inst_35.INIT_RAM_03 = 288'h9A45229138A44E27138A45229149A4D269349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_04 = 288'hAA552A954AA552A9549A5526934AA4D26954AA4D26934AA4D269549A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_05 = 288'hAA552E974AA552A954AA552A954AA5D2A954AA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_35.INIT_RAM_06 = 288'hE3F1F8FA6B2A890482412080544B1D92C964A1D92894381D8943AE54B1A6954AA552A954;
defparam promx9_inst_35.INIT_RAM_07 = 288'h11395CAE461A8904E20379E428130A0904614098A8840A298504E392D164B66C369B4DA6;
defparam promx9_inst_35.INIT_RAM_08 = 288'h9A4D2291389C4E271389C4E271379BCDE6D3692C964B158A44A00FE6DB256A832A1003A0;
defparam promx9_inst_35.INIT_RAM_09 = 288'h9A4D269349A4D229349A4D269348A4D269149A45269349A4D269349A45229348A4526934;
defparam promx9_inst_35.INIT_RAM_0A = 288'h6934DE6F389C4DE6D2591C4D24140D34609169BCE27138A45229149A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_0B = 288'h9A4D269349A4D267139A4D267349A4CE693489CCE693389C4E271389C4DE6F36934964D2;
defparam promx9_inst_35.INIT_RAM_0C = 288'h9A4D269348A452673499C5269148A4D269349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_0D = 288'hAA552A9549A552A9549A5526934AA5526954AA4D2A954AA4D269549A4D2A9349A4D26934;
defparam promx9_inst_35.INIT_RAM_0E = 288'hAA552A954AA552A954AA552A954AA552A954AA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_35.INIT_RAM_0F = 288'hC361B4DA7D3F1F8F86B2B0C82A2510030B63B2592C964B25928944A1C0E0663B0A962954;
defparam promx9_inst_35.INIT_RAM_10 = 288'hA5AA4CC6400F8506E47231186A240C8FCDC850188C28241208C2C2B1410C282724920986;
defparam promx9_inst_35.INIT_RAM_11 = 288'h8A4D269348A4D2291489C52271389C4E26F379BCDE6F369BC9A4D2692C962912803FDDAD;
defparam promx9_inst_35.INIT_RAM_12 = 288'h9A4D269348A45269349A4D269349A45269349A4D229348A45229149A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_13 = 288'h79BCDE6F379C4E271389BCDE6F2588C0826161EB8A0B269BCE271389C5269349A4D26914;
defparam promx9_inst_35.INIT_RAM_14 = 288'h99CCE69349A4CE693499CCE69349A4D2673399CCE69339A4CE271389C4E271389C4E2713;
defparam promx9_inst_35.INIT_RAM_15 = 288'h9A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D26933;
defparam promx9_inst_35.INIT_RAM_16 = 288'hAA552A954AA5526954AA552A9549A55269349A4D269349A4D269549A552A9549A4D26934;
defparam promx9_inst_35.INIT_RAM_17 = 288'h922122934AA552A954AA552A954AA552A954AA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_35.INIT_RAM_18 = 288'h4138E8B45C369F4DA7E3F1F8F86A2A0904823108A8764B2592C964B2512874491C0A4703;
defparam promx9_inst_35.INIT_RAM_19 = 288'h58A44E03007F3AD8C942993C3E172B9588C351A890303E2C994282409850463611118A81;
defparam promx9_inst_35.INIT_RAM_1A = 288'h9A45269349A44E69349A452291489C52271389C4E26F379BCE26F379BCDE6F369349A4B2;
defparam promx9_inst_35.INIT_RAM_1B = 288'h9A4D227148A4D229149A4D269349A45269349A4D269148A4D229149A45229148A44E6934;
defparam promx9_inst_35.INIT_RAM_1C = 288'h89C4E271389BCDE71389C4E271389BCDE6F259140C241B283D24D379C4E271389C522914;
defparam promx9_inst_35.INIT_RAM_1D = 288'h9A4CE69349A4D2693399CD2673489CCE673499CCE673399CCE273399C4E271389CCE2713;
defparam promx9_inst_35.INIT_RAM_1E = 288'h9A4D269349A4D269349A4D269349A4D267349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_1F = 288'hAA552A954AA5526954AA4D26934AA552A934AA4D269349A4D269349A55269349A4D26934;
defparam promx9_inst_35.INIT_RAM_20 = 288'hA248E07038239A69349A552A954AA552A954AA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_35.INIT_RAM_21 = 288'h41590464330A0A4965A2D9B0DA6E3F1F4D8661985048200612C964B2592C964B2592C943;
defparam promx9_inst_35.INIT_RAM_22 = 288'h79BCDE6D26934962B1381401FCEA62A50C63F0005CAE46239146A240C0F4803412090461;
defparam promx9_inst_35.INIT_RAM_23 = 288'h9A4D229148A45229149A45229148A45269148A452291389C4E271389C4E271389BCE26F3;
defparam promx9_inst_35.INIT_RAM_24 = 288'h89C4E27138A45227148A45269349A4D269148A452291399C4E671389CD267339A44E2914;
defparam promx9_inst_35.INIT_RAM_25 = 288'h89C4E271389C4E271389C4E271389C4E271389C4DE6F3692C41F8D07AC9A4F379C4E2713;
defparam promx9_inst_35.INIT_RAM_26 = 288'h9A4D269349A4D267339A4D2693499CCE673389CCE671389C4E271389C4E673389C4E2713;
defparam promx9_inst_35.INIT_RAM_27 = 288'h9A4D269349A4D269349A4D269349A4D269349A4D269349A4D2673499CD269349A4D26934;
defparam promx9_inst_35.INIT_RAM_28 = 288'hAA552A954AA552A954AA55269349A4D2A954AA552A9549A4D269549A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_29 = 288'hB2592C964A248E06C240F2E27349A552A954AA552A954AA552A954AA552A954AA552A954;
defparam promx9_inst_35.INIT_RAM_2A = 288'hD2790C482311854443A01050524A2D168BA7E3E9F4D6541184C440B2D92C964C25930964;
defparam promx9_inst_35.INIT_RAM_2B = 288'h89C4E271379BCE26F379349A4D259244E27017F3E98A84298BC04272391C8C451A098503;
defparam promx9_inst_35.INIT_RAM_2C = 288'h89C4E27148A452273489C4E69148A4D229148A45229139A452691389C4E271389C4E2713;
defparam promx9_inst_35.INIT_RAM_2D = 288'h89C4E27138A452271489C4E271389C4E29148A452291489CD2293389C4E271389CD22713;
defparam promx9_inst_35.INIT_RAM_2E = 288'h89C4E271389C4E271389C4E271389BCE26F389C4E271389C4E26F3793CDA4B269349E713;
defparam promx9_inst_35.INIT_RAM_2F = 288'h9A4D2693399CD269339A4D227139A4D2271389C4E673489CCE273389C4E671389C4E6713;
defparam promx9_inst_35.INIT_RAM_30 = 288'h9A4D269349A4D269349A4D269349A4D269349A4D269349A4D2693399CD267349A4D26933;
defparam promx9_inst_35.INIT_RAM_31 = 288'hAA552A934AA552A954AA4D2A9549A4D269349A4D2A9349A4D2A9549A55269549A4D26934;
defparam promx9_inst_35.INIT_RAM_32 = 288'hB2592C964B25928743A248E072351346273499CD26954AA4D2A954AA552A934AA5526954;
defparam promx9_inst_35.INIT_RAM_33 = 288'h7230D46A25148F0CA020985468062A00C282B2D9ACB86D361ACB0441208C223A1E0EC964;
defparam promx9_inst_35.INIT_RAM_34 = 288'h89C4E671389CCE271389C4E271389BCDE4F279349A4B2489405FCEA5A210A4200B11C8C4;
defparam promx9_inst_35.INIT_RAM_35 = 288'h89C4E271389C4E29148A452273489C5227138A452271389C4E27148A452271389C4E2713;
defparam promx9_inst_35.INIT_RAM_36 = 288'h79C4DE71389C4E271389C4E271389C4E271389C4E27138A45227138A452273399C4E2713;
defparam promx9_inst_35.INIT_RAM_37 = 288'h89C4E271389C4E271399C4E271389C4E271389C4E271389C4E271389C4E271389BCDE6F3;
defparam promx9_inst_35.INIT_RAM_38 = 288'h9A4D269339A4D269339A4CE691399CCE273489CCE271389C4E273389C4E271389C4E2713;
defparam promx9_inst_35.INIT_RAM_39 = 288'h9A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D2693399CCE6734;
defparam promx9_inst_35.INIT_RAM_3A = 288'h9A4D26954AA552A954AA552A954AA552A934AA4D2A9549A4D269349A4D269349A4D26934;
defparam promx9_inst_35.INIT_RAM_3B = 288'hB2592C964B2592C964B25928744A24924744413CA27339A4D269349A552A954AA4D26934;
defparam promx9_inst_35.INIT_RAM_3C = 288'h5308402C47239186C351208832372D1082C220418806151516CB45B2D95C6824118A4164;
defparam promx9_inst_35.INIT_RAM_3D = 288'h89C4E273389C4E271389C4E271389C4E271389C4DE6F379BC9A4D2592C5225017F3A1687;
defparam promx9_inst_35.INIT_RAM_3E = 288'h89C4E271389C4E271389C4E271389C4E271389C4E271389C4E291399CCE271389C4E2713;
defparam promx9_inst_35.INIT_RAM_3F = 288'h89C4E271389C4E271389C4DE71389C4E271389C4E271389C4E271389C4E271389C4E2713;

pROMX9 promx9_inst_36 (
    .DO({promx9_inst_36_dout_w[26:0],promx9_inst_36_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_47),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_36.READ_MODE = 1'b1;
defparam promx9_inst_36.BIT_WIDTH = 9;
defparam promx9_inst_36.RESET_MODE = "SYNC";
defparam promx9_inst_36.INIT_RAM_00 = 288'h89C4E271389C4E271389C4E271399C4E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_01 = 288'h9A4D2693499CD2673499CCE67339A4D2671389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_02 = 288'h9A55269349A45269349A4D269348A4D269349A4D269149A4D269349A4D269148A4D26934;
defparam promx9_inst_36.INIT_RAM_03 = 288'hAA552A9549A552A934AA552A9549A5526954AA4D2A9349A4D2A9549A4D269349A4D26934;
defparam promx9_inst_36.INIT_RAM_04 = 288'h205018543B1D92C964B2592C964B250E8944A2491C4E3633CE271399CD269349A4D26934;
defparam promx9_inst_36.INIT_RAM_05 = 288'h489405FCE85219482210B91C8E461B0D4642F09854482511868C404128A4904512090482;
defparam promx9_inst_36.INIT_RAM_06 = 288'h89C4E271389C4E271389C4E671399CCE671389C4E271389C4E271389BCDE6F269349A4B1;
defparam promx9_inst_36.INIT_RAM_07 = 288'h89C4E271389C4E271389C4E271389C4E271389C4E271389C4E271389C4E271399C4E2733;
defparam promx9_inst_36.INIT_RAM_08 = 288'h89C4E271389C4E271379C4E271389C4E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_09 = 288'h89C4E271389C4E271389C4E271389C4E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_0A = 288'h9A4D267349A44E69349A4CE673499CD2673399CCE271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_0B = 288'h9A4D269349A4D269349A4D229349A4D269349A4D269349A4D269349A45229349A4D26914;
defparam promx9_inst_36.INIT_RAM_0C = 288'hAA4D26934AA4D2A954AA4D269349A4D2A934AA4D269349A4D269349A55269349A4D26934;
defparam promx9_inst_36.INIT_RAM_0D = 288'h40A0442C0B2D0E86E2B258EC964B25928764A1D0E8AE09240E46C368BCE271399CD26934;
defparam promx9_inst_36.INIT_RAM_0E = 288'h79BCDE4D258AC4E05007635D28652084C4E47239186A341985048251388830320984C482;
defparam promx9_inst_36.INIT_RAM_0F = 288'h89C4E271389C4E671389C4E271399C4E271399C4E271389C4E271389C4E271389C4E26F3;
defparam promx9_inst_36.INIT_RAM_10 = 288'h89C4E271389C4DE71389C4E271389C4E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_11 = 288'h89C4E271389C4E271389C4DE71389C4E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_12 = 288'h89C4E271379C4E271389C4E271389C4E271389BCE271389C4E271389C4DE71389BCDE713;
defparam promx9_inst_36.INIT_RAM_13 = 288'h9A4CE673499CD2693489C4E273399CCE273399CCE673389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_14 = 288'h9A4D267349A4D269349A4D2693499CD2273399CCE67349A4D269339A4D269339A4D26934;
defparam promx9_inst_36.INIT_RAM_15 = 288'h99CD269349A4D269349A4D269349A4D269349A55269349A4D269349A4D269349A4D26934;
defparam promx9_inst_36.INIT_RAM_16 = 288'h6218484201018B4943A158EC74370D12C964B25928764A1D128900F0C8E46C6793CE2713;
defparam promx9_inst_36.INIT_RAM_17 = 288'h89C4E271389C4DE6F269349629138143DF6D74995084151B9588C490C1D422261090C180;
defparam promx9_inst_36.INIT_RAM_18 = 288'h89C4E271389C4E271389C4E271389C4E271389C4E691399C4E27139A44E273489C4E2713;
defparam promx9_inst_36.INIT_RAM_19 = 288'h89BCE271389C4E271389C4E26F389C4E271389C4DE71389C4DE71389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_1A = 288'h89BCE271389BCDE6F379C4E271389C4E271389C4E271389C4E271389BCDE71389C4E2713;
defparam promx9_inst_36.INIT_RAM_1B = 288'h89C4E271389C4E271389C4DE71389BCE271379BCDE71389C4E271389C4E271389BCDE713;
defparam promx9_inst_36.INIT_RAM_1C = 288'h99C4E673389C4E671399C4E271399C4E27339A4D267339A4CE691399C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_1D = 288'h9A4D269349A4D269139A4D2693399CCE671399C4E673499CD2271399CCE27339A44E6933;
defparam promx9_inst_36.INIT_RAM_1E = 288'h7944E271389CD269349A4D26934AA4D2A9349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_36.INIT_RAM_1F = 288'h30A0584E25128F4BC5D2E12C763B1D8EC763B238AC964B25928743A1D92872391C8D446F;
defparam promx9_inst_36.INIT_RAM_20 = 288'h89C4E271389C4E271389C4DE6F3693C9A4B258A40A02FF75B1D26542005C8E562A9148A2;
defparam promx9_inst_36.INIT_RAM_21 = 288'h89C4E271389C4E271389C4E271389C4E271389C4E271389CCE271389C4E271389C4E6913;
defparam promx9_inst_36.INIT_RAM_22 = 288'h89C4E26F379C4E271389BCE26F379C4E271389C4E271379BCDE6F379C4E271389C4DE713;
defparam promx9_inst_36.INIT_RAM_23 = 288'h89C4E26F389BCDE71379BCDE6F379BCE271389C4DE6F389C4E26F379BCDE6F389C4E26F3;
defparam promx9_inst_36.INIT_RAM_24 = 288'h89C4E271389C4E26F379C4E26F379BCDE6F389C4E26F389BCDE71389BCE26F389BCE2713;
defparam promx9_inst_36.INIT_RAM_25 = 288'h89CCE671389C4E67139A44E671389CCE671389C4E273399CCE271389C4E273389C4E2713;
defparam promx9_inst_36.INIT_RAM_26 = 288'h9A4D269349A4D2693499C4E271389C4E271389CD2673389CCE273389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_27 = 288'h81C0D06D279BCE271389C4E69349A4D269349A4D269349A4D269349A4D269349A4D26934;
defparam promx9_inst_36.INIT_RAM_28 = 288'h62B1548A26118902C250E0FCDC5D26130983B1D8EC763B250DC564B2592C964A1D0E8723;
defparam promx9_inst_36.INIT_RAM_29 = 288'h89C4E273489C4E69139A44E271389C4E271379BCDE4D2692C52270280BF9D6C75218C863;
defparam promx9_inst_36.INIT_RAM_2A = 288'h79C4DE71379BCE271379BCE271389BCE271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_2B = 288'h89C4DE6F379BCDE71389C4DE71389BCDE71379BCDE71379C4E271379C4DE71379C4DE713;
defparam promx9_inst_36.INIT_RAM_2C = 288'h79BCDE6F379C4DE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F389BCE26F379BCDE713;
defparam promx9_inst_36.INIT_RAM_2D = 288'h89C4E271389BCDE71389BCE26F389BCDE6F379BCDE6F379BCDE6F379C4DE6F379BCDE6F3;
defparam promx9_inst_36.INIT_RAM_2E = 288'h89C4E271389C4E271389C4E673389C4E271389C4E271389C4E273389CCE271389C4E2713;
defparam promx9_inst_36.INIT_RAM_2F = 288'h9A4D2693499C4E693489CD269349A44E271389C4E273389CCE271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_30 = 288'hB250E8723A2184DCF379C4E271389CD2673399CD2693499CD269349A4D269349A4D26934;
defparam promx9_inst_36.INIT_RAM_31 = 288'hD75B214A813F99D460F1B0DC6822030BC9C5D26130963B1D8EC763B1D0EC902A1D0E8743;
defparam promx9_inst_36.INIT_RAM_32 = 288'h89C4E273489CCE69139A4D269349A44E273399CCE271389C4DE6F2793C9A2B1489C0A1EF;
defparam promx9_inst_36.INIT_RAM_33 = 288'h79BCDE6F379BCDE71379BCDE6F379BCE271379C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_34 = 288'h89BCE271379C4DE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379C4E271379BCDE6F3;
defparam promx9_inst_36.INIT_RAM_35 = 288'h79BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE71389BCE271379BCDE713;
defparam promx9_inst_36.INIT_RAM_36 = 288'h89C4E271389C4E271379BCDE71379BCDE6F379BCDE6F379BCDE6F379BCDE6F379C4DE6F3;
defparam promx9_inst_36.INIT_RAM_37 = 288'h89C4E271389C4E271389C4E271389C4E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_38 = 288'h9A4D2273499CD2693499CD2673499C4E271389C4E271389C4E273389C4E271389C4E2713;
defparam promx9_inst_36.INIT_RAM_39 = 288'h9250E8743A1D0E46E261295A4D279C4E271389CCE69349A4D269349A4D269349A4D26934;
defparam promx9_inst_36.INIT_RAM_3A = 288'h692C5227017FBF5D4C85AA85104B2B0D50853090102C1C260F0783B1D8EC783B2512C824;
defparam promx9_inst_36.INIT_RAM_3B = 288'h89C4E271389C4E271389C4E69139A4D2271399CCE673389CCE671389C4E26F379BC9A4D2;
defparam promx9_inst_36.INIT_RAM_3C = 288'h79BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCE26F379C4E2713;
defparam promx9_inst_36.INIT_RAM_3D = 288'h79BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379C4DE6F379BCDE6F3;
defparam promx9_inst_36.INIT_RAM_3E = 288'h79C4DE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F3;
defparam promx9_inst_36.INIT_RAM_3F = 288'h89C4E271389C4E271389C4E271379C4DE6F379BCDE6F379BCDE6F379BCDE4F379BCDE6F3;

pROMX9 promx9_inst_37 (
    .DO({promx9_inst_37_dout_w[26:0],promx9_inst_37_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_49),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_37.READ_MODE = 1'b1;
defparam promx9_inst_37.BIT_WIDTH = 9;
defparam promx9_inst_37.RESET_MODE = "SYNC";
defparam promx9_inst_37.INIT_RAM_00 = 288'h89C4E26F389C4E271389C4E271389C4E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_37.INIT_RAM_01 = 288'h99CCE27349A4D2693399CD267339A44E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_37.INIT_RAM_02 = 288'hA1A12461095D164722A1C8DC544312C5A2F389C4E271389CD269349A44E27139A4D22733;
defparam promx9_inst_37.INIT_RAM_03 = 288'h89C4DE4F27934962B1389401FEED75B658A93128BD02120280826150C0A8743B1D8EC744;
defparam promx9_inst_37.INIT_RAM_04 = 288'h89C4DE6F389C4E271389C4E271389C4E69139A4D2271389CCE673399CCE673399C4E2713;
defparam promx9_inst_37.INIT_RAM_05 = 288'h79BCDE4F379BCDE6F379BC9E6F279BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE713;
defparam promx9_inst_37.INIT_RAM_06 = 288'h79BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F3793CDE4F379BCDE6F379BCDE6F3;
defparam promx9_inst_37.INIT_RAM_07 = 288'h79BCDE4F3793C9E4F379BC9E4F3793CDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F3;
defparam promx9_inst_37.INIT_RAM_08 = 288'h89C4E271389C4E271389BCE271379C4DE6F379BCDE6F379BCDE6F379BCDA4F379BCDE6F3;
defparam promx9_inst_37.INIT_RAM_09 = 288'h89C4E271389C4E271389C4E271389C4E271389BCE271389C4E271389C4E271379C4E2713;
defparam promx9_inst_37.INIT_RAM_0A = 288'h99CCE673399CCE671399CCE27339A4D2693399CCE273389CCE26F379C4E271379C4E2713;
defparam promx9_inst_37.INIT_RAM_0B = 288'hA1592C724B1E1BDE10F7B26492491C0E8881173C9E51289C4E271389CCE691389CD26733;
defparam promx9_inst_37.INIT_RAM_0C = 288'h89C4E671389C4E271379BC9A4D258A44A03017FBB9D8DA61229A2803B8C0FAA51285C303;
defparam promx9_inst_37.INIT_RAM_0D = 288'h79BC9E713793CDE6F379C4E271389C4E271389C4E273399CCE273399CCE673399CCE6733;
defparam promx9_inst_37.INIT_RAM_0E = 288'h79BC9E6F2793C9A4F379BC9E4F279BCDE4D279BC9E6F279BCDE6F379B49A4F379BCDE6F3;
defparam promx9_inst_37.INIT_RAM_0F = 288'h79BCDE4F379BCDE6F379BCDE4F379BCDE4F379BC9E6F279BCDE4F3793C9E4F379BCDE4F3;
defparam promx9_inst_37.INIT_RAM_10 = 288'h79BCDE6D2693CDE4D2793C9E6F2793C9E4F2693C9E4F279BCDE6F379BC9E6F379BC9E6F3;
defparam promx9_inst_37.INIT_RAM_11 = 288'h89C4DE71389C4E271389C4E271389BCDE71379BCDE6F379BCDE6F379BC9A4D2693C9E6F3;
defparam promx9_inst_37.INIT_RAM_12 = 288'h79C4E271389C4E271389C4E271379C4E271389C4E271389C4E271389C4E26F389C4E2713;
defparam promx9_inst_37.INIT_RAM_13 = 288'h99CCE671399CCE673499CD2671399CCE67349A44E673389C4E271389C4E271389C4DE6F3;
defparam promx9_inst_37.INIT_RAM_14 = 288'h24192CC8C82C848745F77BFDFCFE7F388F0381C8D84C768B49E51289C4E271389C4E6713;
defparam promx9_inst_37.INIT_RAM_15 = 288'h99CCE673399CCE671389C4E271389BCDE6D2692C964913814061EFE7E365848209045021;
defparam promx9_inst_37.INIT_RAM_16 = 288'h79BCDE6F2793C9E6F279BCDE6F389BCDE71389C4E271389C4E271399CCE671399CCE6733;
defparam promx9_inst_37.INIT_RAM_17 = 288'h79349E6F379349A4F279349E4F2693C9A4D269349A4F279349E4F3693CDE6D2693CDE6F3;
defparam promx9_inst_37.INIT_RAM_18 = 288'h79BCDE6F2793CDE4F2793C9E4F2793C9E4F3793C9E6F2793CDE4F279349E6F279349E4F3;
defparam promx9_inst_37.INIT_RAM_19 = 288'h69349A4D279349A4F269349E4D269349E4D279349A4D269349A4D2693CDA4F369349E4F3;
defparam promx9_inst_37.INIT_RAM_1A = 288'h79C4E271379BCE26F379C4DE6F389C4E271389BCDE6F379BCDE6F379BC9E4F2793C9A4D2;
defparam promx9_inst_37.INIT_RAM_1B = 288'h79C4DE51379BCDE6F379BCE271389C4E26F379BCDE6F389C4DE6F379C4DE71389C4DE713;
defparam promx9_inst_37.INIT_RAM_1C = 288'h89C4E271389CCE271389CCE27339A44E693489C4E273499C4E271389CCE671389C4DE713;
defparam promx9_inst_37.INIT_RAM_1D = 288'h85A255469C2D9704E5358D59B2350D975DCED7EBB1BC48230A50B179349E71389C4E2713;
defparam promx9_inst_37.INIT_RAM_1E = 288'h99CCE67349A4CE67339A4D2673399CCE671389C4E26F379BC9A4D258A44E050187BF9D6D;
defparam promx9_inst_37.INIT_RAM_1F = 288'h69349E4F3693C9E4F379BC9E4F2793CDE6F379C4DE51379C4DE71379BCE271389C4E6733;
defparam promx9_inst_37.INIT_RAM_20 = 288'h693C9A4D269349A4F2693C9E4F269349A4D2693C9A4D269349A4F369349A4D269349A4F3;
defparam promx9_inst_37.INIT_RAM_21 = 288'h793C9E4D2693C9A4F2793C9E6F2793C9E4F279BCDA4F369349A4D269349E4F279B49A4D2;
defparam promx9_inst_37.INIT_RAM_22 = 288'h693CDA4D2793CDA4D279B49A4D269349A4D2693CDA4D279349A4D269349E4F2693C9E4D2;
defparam promx9_inst_37.INIT_RAM_23 = 288'h79C4E26F379C4DE6F379BCDE6F379BCDE6F379BCDE6F379BCDE6F379BCDE4F279349A4D2;
defparam promx9_inst_37.INIT_RAM_24 = 288'h89C4E271389BCDE4F379BCDE6F379BCDE6F379BCDE6F389BCE26F379C4DE71379BCDE6F3;
defparam promx9_inst_37.INIT_RAM_25 = 288'h89C4E271389C4E271399CCE271399C4E691389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_37.INIT_RAM_26 = 288'h38940A00FD75B658A94491FCA0372D1F926A04E17C68295DB6160471B9962D1793C9E713;
defparam promx9_inst_37.INIT_RAM_27 = 288'h89C4E271389C4E673499CCE67339A4CE673399CCE273389C4E271389C4DE6D2693496491;
defparam promx9_inst_37.INIT_RAM_28 = 288'h69349A4D2693CDA4D2693C9A4D2793C9E4F379B49E6F279BCDE71379C4E271389C4E2713;
defparam promx9_inst_37.INIT_RAM_29 = 288'h79B49A4D2693C9A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D2;
defparam promx9_inst_37.INIT_RAM_2A = 288'h69349A4D279349A4D2793CDE6D269349A4D269349E4F269349E4D279B49A4D269349A4F2;
defparam promx9_inst_37.INIT_RAM_2B = 288'h69349E4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D279B49A4D2;
defparam promx9_inst_37.INIT_RAM_2C = 288'h79BCDE6F279BCDE6F279BC9E4F3793CDE6F379BCDE6F389BCDE6F379BCDA4F279BCDA4D2;
defparam promx9_inst_37.INIT_RAM_2D = 288'h89C4E271389C4E26F379BCDE4D279BCDE6F379BCE26F379BCDE6F379BCE26F379BCDE6F2;
defparam promx9_inst_37.INIT_RAM_2E = 288'h7944E271389C4E271389CCE671389C4E271389C4E271389C4E271389C4E271389C4E2713;
defparam promx9_inst_37.INIT_RAM_2F = 288'h79BCDA6B2592C922501803F5D8DB642D90E793CA24F48B46A2CD4662D854CC3C52C9A2F2;
defparam promx9_inst_37.INIT_RAM_30 = 288'h89C4E271389CCE271389CCE273399CCE673399CCE673399CCE673399C4E671389C4DE6F3;
defparam promx9_inst_37.INIT_RAM_31 = 288'h69349A4D269349A4D269349A4D269349A4D2693C9A4D269349E4F2793CDE6F379C4E26F3;
defparam promx9_inst_37.INIT_RAM_32 = 288'h69349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D2;
defparam promx9_inst_37.INIT_RAM_33 = 288'h69349A4D269349A4D269349A4D269349A4D269349A4D269349A4D279349A4D269349A4D2;
defparam promx9_inst_37.INIT_RAM_34 = 288'h693CDE4D269349A4D269349A4D269349A4D2692C9A4D269349A4D269349A4D26934964D2;
defparam promx9_inst_37.INIT_RAM_35 = 288'h79BCDE6F379BCDE6F379BC9E6F3693CDE6F379BC9E6F379BCDE6F379BCDA4F279BC9E4F2;
defparam promx9_inst_37.INIT_RAM_36 = 288'h89C4E271389C4E271379C4E26F379BCDE4F279BCDA4F379BCDE6F379BCDE6F379BC9E6F3;
defparam promx9_inst_37.INIT_RAM_37 = 288'h58B49A4D279BCE271389C4E271389CCE271389C4E271389C4E671389C4E271389C4E2713;
defparam promx9_inst_37.INIT_RAM_38 = 288'h89C4E271389C4DE6F369B4964B248A44A05007FBB9B6BA54A65349A45A61129A4D245C8F;
defparam promx9_inst_37.INIT_RAM_39 = 288'h793CE271389C4E271389C4E271389C4E671399CCE673399CCE67339A4D2673399CCE2713;
defparam promx9_inst_37.INIT_RAM_3A = 288'h6934964B269349A4D26934964D269349A4B269349A4D269349A4D279349A4F2793C9E4F2;
defparam promx9_inst_37.INIT_RAM_3B = 288'h69349A4D269349A4D269349A4D2692C9A4D259349A4D269349A4D269349A4B259349A4B2;
defparam promx9_inst_37.INIT_RAM_3C = 288'h69349A4D2692C9A4B269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D2;
defparam promx9_inst_37.INIT_RAM_3D = 288'h69349A4D269349A4D269349A4D269349A4D269349A4D2692C964D269349A4D259349A4D2;
defparam promx9_inst_37.INIT_RAM_3E = 288'h79BCDE4F2793CDE6F379BCDE4F379BC9A4D269349A4D269349E6F3793C9E6F2793C9E4F3;
defparam promx9_inst_37.INIT_RAM_3F = 288'h89C4DE71379C4E271379C4E26F379BCDE4F3793C9E6F269349E6F369349E6D279BCDE4F2;

pROM prom_inst_38 (
    .DO({prom_inst_38_dout_w[30:0],prom_inst_38_dout[9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_38.READ_MODE = 1'b1;
defparam prom_inst_38.BIT_WIDTH = 1;
defparam prom_inst_38.RESET_MODE = "SYNC";
defparam prom_inst_38.INIT_RAM_00 = 256'h000000000000000200000000000F3C000FF98000000020000000000000000033;
defparam prom_inst_38.INIT_RAM_01 = 256'h00000000100000000003DFC001FF1000000006000200000000000005FFFFF000;
defparam prom_inst_38.INIT_RAM_02 = 256'h000000000001C5FE007FE300000000400000000000000000BFFFFFC000000000;
defparam prom_inst_38.INIT_RAM_03 = 256'h0000309FFC1FFC600000000400000000000000001BFFFFFF0000000000000000;
defparam prom_inst_38.INIT_RAM_04 = 256'hFFFFFF0C000000004000000000000000037FFFFFF80000000000000000020000;
defparam prom_inst_38.INIT_RAM_05 = 256'h800000000C00000000000000006FFF9FFEE00000000000000000081000000E77;
defparam prom_inst_38.INIT_RAM_06 = 256'h00C00000000000000005FFF0FFF780000000000000000000000003CE3FFFFFE1;
defparam prom_inst_38.INIT_RAM_07 = 256'h000000000000BFFE03FF1E0000000000000000000000007FC3FFFFFC70000000;
defparam prom_inst_38.INIT_RAM_08 = 256'h00001BFFC00FF07000000000000000000000000FF03FFBFF8E00000000080000;
defparam prom_inst_38.INIT_RAM_09 = 256'hFC003F81C00000000000000000000001FF13FF7FF9C0000000008000C0000000;
defparam prom_inst_38.INIT_RAM_0A = 256'h0700000000000000000000003FC01FF3EF9C000000001800000000000000037F;
defparam prom_inst_38.INIT_RAM_0B = 256'h000000000000000003F0007F86FB800000000180000000000000002FFF8000FC;
defparam prom_inst_38.INIT_RAM_0C = 256'h00000000001E1009E00FB800000000100000000000000002FFF00003F04C0000;
defparam prom_inst_38.INIT_RAM_0D = 256'h0000C7001200FB80000000010001000000000000C7FE00000FC0600000000000;
defparam prom_inst_38.INIT_RAM_0E = 256'h00400F98000000001000000000000000047FA000007F83800000000000000000;
defparam prom_inst_38.INIT_RAM_0F = 256'h800000000300000000000000018FFC000007FC4E0000000000000000000100F0;
defparam prom_inst_38.INIT_RAM_10 = 256'h00300000000000000008FF8000007FF730000000000000000000003E000000F9;
defparam prom_inst_38.INIT_RAM_11 = 256'h0000000000031FFF00000FFFDCC000000000000000000000E0020007B0000000;
defparam prom_inst_38.INIT_RAM_12 = 256'h000033FFFC0001FFFF730000000000000000000000003E007B00000000020001;
defparam prom_inst_38.INIT_RAM_13 = 256'hFFF0001FFFFD8C600000000000000000000001E0033000000000200000000000;
defparam prom_inst_38.INIT_RAM_14 = 256'hFFFFFA60000000000000000010000004001300000000020000000000000003FF;
defparam prom_inst_38.INIT_RAM_15 = 256'h0000000000000000010000000000300000000020002000000000003FEFFFC003;
defparam prom_inst_38.INIT_RAM_16 = 256'h000000000000000000000700000000060000000000000003FFFF7D806FFFFFF0;
defparam prom_inst_38.INIT_RAM_17 = 256'h00008000000000600000000040000000000000003FFFFEE600B2BFF8E0000000;
defparam prom_inst_38.INIT_RAM_18 = 256'h0000010E00000000040004000000000003FFFFFFF80C00FF818C000000000000;
defparam prom_inst_38.INIT_RAM_19 = 256'hC000000000C0000000000000001FFFFFFEF04007F803F0000000000000000400;
defparam prom_inst_38.INIT_RAM_1A = 256'h000C0000000000000000F3FFFFFFE8003F0007C00000000000000020000000D0;
defparam prom_inst_38.INIT_RAM_1B = 256'h8000000000000F8FFFF9F70003F0003F00000000000000010180001C18000000;
defparam prom_inst_38.INIT_RAM_1C = 256'h0000007C3FF807C0003E0001F800000000000000041FC00D0300000000008000;
defparam prom_inst_38.INIT_RAM_1D = 256'hCAFF001F0001E0001FC000000000000000107DE7007000000000000000000000;
defparam prom_inst_38.INIT_RAM_1E = 256'h7E003C0000FE0000000000000000601E400C0000000002000200000000000003;
defparam prom_inst_38.INIT_RAM_1F = 256'h000FF00000000000000001C0000380000000000400100000000000000E07F800;
defparam prom_inst_38.INIT_RAM_20 = 256'h0000000000000002F000E000000000004004000000000000007CFFE000F007C0;
defparam prom_inst_38.INIT_RAM_21 = 256'h000000000E2078000000000004002000000000000001F9FF800380780000FF80;
defparam prom_inst_38.INIT_RAM_22 = 256'h000FFC000000000000C0020000000000000007FFFE000E0F00000FF400000000;
defparam prom_inst_38.INIT_RAM_23 = 256'h00000000000C0120000000000000001F7FF80038E00000FEA000000000000000;
defparam prom_inst_38.INIT_RAM_24 = 256'h000880120000000000000000FDFFC001FC00000FEE0000000000000000000000;
defparam prom_inst_38.INIT_RAM_25 = 256'h200000000000000003EFFF0007800000FEF00000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_26 = 256'h00000000000FFFFA003000001FFF800000000000000000000000000000001000;
defparam prom_inst_38.INIT_RAM_27 = 256'h00003FFFD801000001FE38000000000000000000000000000000060002000000;
defparam prom_inst_38.INIT_RAM_28 = 256'hFF400800003FF9C0000000000000000000000000000000000260000000000000;
defparam prom_inst_38.INIT_RAM_29 = 256'h0003FFF4000000000000000000000000000000000024000000000000000000FE;
defparam prom_inst_38.INIT_RAM_2A = 256'hC0000000000000000000000000000000000040000000000000000003FBFF0040;
defparam prom_inst_38.INIT_RAM_2B = 256'h00000000000000000000000000000000000000000000000007CFFC0600007FFF;
defparam prom_inst_38.INIT_RAM_2C = 256'h0000000000000000000001000000000000000000001F7FF0300007FFFC000000;
defparam prom_inst_38.INIT_RAM_2D = 256'h0000000000000000000000000000000000007DFF810000FFFFC0000000000000;
defparam prom_inst_38.INIT_RAM_2E = 256'h000000000000000000000000000001FFFE08001FFFF800000000000000000000;
defparam prom_inst_38.INIT_RAM_2F = 256'h000000000000000000000007FFF84001FFFF8000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_30 = 256'h00000000000000001FFF02003FFFF80000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_31 = 256'h00000000007FF8100FFFEF000000000000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_32 = 256'h0003FF5C87FFFE70000000000000000000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_33 = 256'hFFFFFFFE00000000000000000000000000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_34 = 256'hE000000000000000000000000000000000000000000000000000000000000FFF;
defparam prom_inst_38.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000003FFFFFFFFF;
defparam prom_inst_38.INIT_RAM_36 = 256'h000000000000000000000000000000000000000000000001FA7FFFFFFC000000;
defparam prom_inst_38.INIT_RAM_37 = 256'h000000000000000000000000000000000000000007E3FFFFFFC0000000000000;
defparam prom_inst_38.INIT_RAM_38 = 256'h00000000000000000000000000000000001F03FFCFF800000000000000000000;
defparam prom_inst_38.INIT_RAM_39 = 256'h00000000000000000000000000007FBFF2FF0000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_3A = 256'h0000000000000000000001F2EEFFF00000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_3B = 256'h0000000000000007F153EE000000000000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_3C = 256'h000000000FDE4FC0000000000000000000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_3D = 256'h003FFFB800000000000000000000000000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_38.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000007FFC;

pROM prom_inst_39 (
    .DO({prom_inst_39_dout_w[30:0],prom_inst_39_dout[10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_39.READ_MODE = 1'b1;
defparam prom_inst_39.BIT_WIDTH = 1;
defparam prom_inst_39.RESET_MODE = "SYNC";
defparam prom_inst_39.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFC0001FFFFFFF0000000007FFFFFFFDFFFDFFFFFFFFFFFFFC0;
defparam prom_inst_39.INIT_RAM_01 = 256'hFFFFFFFFE0001FFFFFFC200000000FFFFFFFF9FFF9FFFFFFFFFFFFF800000FFF;
defparam prom_inst_39.INIT_RAM_02 = 256'hFF8003FFFFFE3A00000000FFFFFFFFBFFFBFFFFFFFFFFFFF0000003FFFFFFFFF;
defparam prom_inst_39.INIT_RAM_03 = 256'hFFFFCF200000001FFFFFFFFBFFFBFFFFFFFFFFFFE0000000FFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_04 = 256'h00000003FFFFFFFFBFFFBFFFFFFFFFFFFC00000007FFFFFFFFFFFFFFFFFC007F;
defparam prom_inst_39.INIT_RAM_05 = 256'h7FFFFFFFF3FFFBFFFFFFFFFFFF800000001FFFFFFFFFFFFFFFFFF00FFFFFF180;
defparam prom_inst_39.INIT_RAM_06 = 256'hFF3FFFBFFFFFFFFFFFF8000000007FFFFFFFFFFFFFFFFFFFFFFFFC3000000000;
defparam prom_inst_39.INIT_RAM_07 = 256'hFFFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFF80000000000FFFFFFF;
defparam prom_inst_39.INIT_RAM_08 = 256'hFFFFE0000000000FFFFFFFFFFFFFFFFFFFFFFFF00000000001FFFFFFFFF7FFFB;
defparam prom_inst_39.INIT_RAM_09 = 256'h000000003FFFFFFFFFFFFFFFFFFFFFFE00000000003FFFFFFFFF7FFF3FFFFFFF;
defparam prom_inst_39.INIT_RAM_0A = 256'h00FFFFFFFFFFFFFFFFFFFFFFC00000000003FFFFFFFFE7FFF7FFFFFFFFFFFC00;
defparam prom_inst_39.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFF800000000007FFFFFFFFE7FFF7FFFFFFFFFFFC000000000;
defparam prom_inst_39.INIT_RAM_0C = 256'hFFFFFFFFFF000000000007FFFFFFFFEFFFF7FFFFFFFFFFF8000000000003FFFF;
defparam prom_inst_39.INIT_RAM_0D = 256'hFFF000000000007FFFFFFFFEFFFE7FFFFFFFFFFF0000000000001FFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0E = 256'h00000007FFFFFFFFEFFFEFFFFFFFFFFFF00040000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0F = 256'h7FFFFFFFFCFFFEFFFFFFFFFFFE00000000000001FFFFFFFFFFFFFFFFFFFE0000;
defparam prom_inst_39.INIT_RAM_10 = 256'hFFCFFFEFFFFFFFFFFFE00000000000000FFFFFFFFFFFFFFFFFFFE00000000000;
defparam prom_inst_39.INIT_RAM_11 = 256'hFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFFFFFE00000000000FFFFFFF;
defparam prom_inst_39.INIT_RAM_12 = 256'hFFFFC000000000000000FFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFDFFFC;
defparam prom_inst_39.INIT_RAM_13 = 256'h000000000000039FFFFFFFFFFFFFFFFE00000000000FFFFFFFFFDFFFDFFFFFFF;
defparam prom_inst_39.INIT_RAM_14 = 256'h00000019FFFFFFFFFFFFFFFFE00000000000FFFFFFFFFDFFFDFFFFFFFFFFFC00;
defparam prom_inst_39.INIT_RAM_15 = 256'h1FFFFFFFFFFFFFFFFE00000000000FFFFFFFFFDFFF9FFFFFFFFFFFC010000000;
defparam prom_inst_39.INIT_RAM_16 = 256'hFFFFFFFFFFF00000000000FFFFFFFFF9FFFBFFFFFFFFFFFC0000820010000000;
defparam prom_inst_39.INIT_RAM_17 = 256'hFFFF00000000001FFFFFFFFFBFFFBFFFFFFFFFFFC0000118074D400001FFFFFF;
defparam prom_inst_39.INIT_RAM_18 = 256'h00000001FFFFFFFFFBFFF3FFFFFFFFFFFC00000000F3FF000003FFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_19 = 256'h3FFFFFFFFF3FFF7FFFFFFFFFFFE00000010FBFF800000FFFFFFFFFFFFFFFF800;
defparam prom_inst_39.INIT_RAM_1A = 256'hFFF3FFF7FFFFFFFFFFFF0000000017FFC000003FFFFFFFFFFFFFFFC000000000;
defparam prom_inst_39.INIT_RAM_1B = 256'h7FFFFFFFFFFFF000000008FFFC000000FFFFFFFFFFFFFFFE0000000007FFFFFF;
defparam prom_inst_39.INIT_RAM_1C = 256'hFFFFFF800000003FFFC0000007FFFFFFFFFFFFFFF800000000FFFFFFFFFF7FFE;
defparam prom_inst_39.INIT_RAM_1D = 256'h00000000FFFE0000003FFFFFFFFFFFFFFFE00000000FFFFFFFFFE7FFEFFFFFFF;
defparam prom_inst_39.INIT_RAM_1E = 256'h01FFC0000001FFFFFFFFFFFFFFFF80000003FFFFFFFFFC3FFCFFFFFFFFFFFFFC;
defparam prom_inst_39.INIT_RAM_1F = 256'h00000FFFFFFFFFFFFFFFFE0000007FFFFFFFFFC3FFCFFFFFFFFFFFFFF0000000;
defparam prom_inst_39.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFC00001FFFFFFFFFFC3FF9FFFFFFFFFFFFFF800000000FF800;
defparam prom_inst_39.INIT_RAM_21 = 256'hFFFFFFFFF00007FFFFFFFFFFC3FF9FFFFFFFFFFFFFFE000000007F800000007F;
defparam prom_inst_39.INIT_RAM_22 = 256'hFFF003FFFFFFFFFFF83FF1FFFFFFFFFFFFFFF800000001F000000003FFFFFFFF;
defparam prom_inst_39.INIT_RAM_23 = 256'hFFFFFFFFFF83FE1FFFFFFFFFFFFFFFE000000007000000001FFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_24 = 256'hFFF07FE1FFFFFFFFFFFFFFFF000000000000000001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_25 = 256'h1FFFFFFFFFFFFFFFFC00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_26 = 256'hFFFFFFFFFFF000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFE;
defparam prom_inst_39.INIT_RAM_27 = 256'hFFFFC00020000000000047FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFE1FFFFFF;
defparam prom_inst_39.INIT_RAM_28 = 256'h008000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_29 = 256'h00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFF00;
defparam prom_inst_39.INIT_RAM_2A = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFC00000000;
defparam prom_inst_39.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFF800000000000000;
defparam prom_inst_39.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFE000000000000003FFFFFF;
defparam prom_inst_39.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000003FFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFF80000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFE0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_31 = 256'hFFFFFFFFFF800000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_32 = 256'hFFFC00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_33 = 256'h00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_34 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam prom_inst_39.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000;
defparam prom_inst_39.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003FFFFFF;
defparam prom_inst_39.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000003FFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000001007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000100FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFE0010000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFF800E001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3C = 256'hFFFFFFFFF001803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3D = 256'hFFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003;

pROM prom_inst_40 (
    .DO({prom_inst_40_dout_w[30:0],prom_inst_40_dout[11]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_40.READ_MODE = 1'b1;
defparam prom_inst_40.BIT_WIDTH = 1;
defparam prom_inst_40.RESET_MODE = "SYNC";
defparam prom_inst_40.INIT_RAM_00 = 256'h04FFFFFFFFFFFFF61004000000E9A96C004AEF000001B803F3E00000003FF8C4;
defparam prom_inst_40.INIT_RAM_01 = 256'hFFFFFFFDD8004000001DF08B711F20E000001280797E00000003FE1D97EE4C00;
defparam prom_inst_40.INIT_RAM_02 = 256'hFC902E0000071DBA29C1D85E000001200777C00000003FD63516F014007FFFFF;
defparam prom_inst_40.INIT_RAM_03 = 256'h0001BA9FF7F81BF9E000001900F37F0000002FF09E823FC02001FFFFFFFFFF7F;
defparam prom_inst_40.INIT_RAM_04 = 256'hF75F8E8FBE000001500F27F000000DFE3EB40DFF180011FFFFFFFFFFFFC2FE20;
defparam prom_inst_40.INIT_RAM_05 = 256'hD7E000001700E6FE4000007FC67F00D8F878001F3FFFFFFFFDFF9A51000010C7;
defparam prom_inst_40.INIT_RAM_06 = 256'h00401EE7E0000003F8DCF023CB69800177FFFFFFFEFFFE3C000008741FFBE059;
defparam prom_inst_40.INIT_RAM_07 = 256'hFC020013FF1DD701BC2EB28009FFFFFFFFFBFFF8000001816DFEDF0D0A7F0000;
defparam prom_inst_40.INIT_RAM_08 = 256'hFFE392802E8C73200000FFFFFFDBF9FE400000211A4FDBD0184FC800000701E6;
defparam prom_inst_40.INIT_RAM_09 = 256'h27E0313900010DFFF7BE3FFEFC00000F3C0F7CFD1908FC000005B03E2FF40008;
defparam prom_inst_40.INIT_RAM_0A = 256'h6580006FFAF5BB77F7800001ABF693EA0FE31FD100005597E2FFB00367FC35E0;
defparam prom_inst_40.INIT_RAM_0B = 256'hFDE0A40823F8000033FB86E70A7051FEC0000DD47EC7FE8126FFC6AD80FA89CB;
defparam prom_inst_40.INIT_RAM_0C = 256'h1083C000060A08C2E0051D3FF8400085DFFC7FC84FAFF8CDF107B2CC645C0000;
defparam prom_inst_40.INIT_RAM_0D = 256'h01FE446C644181F7FDC0001BDFFC47FF7DFFFF190185FE1A2844C00008C00280;
defparam prom_inst_40.INIT_RAM_0E = 256'h68B0883A7FFE000389FFDDFFEE7FFFE1A044CEFACAE5A9D00000000000000800;
defparam prom_inst_40.INIT_RAM_0F = 256'h27FE7801F81FFB0FFFCFFFFC1B701FC79FA846EC0000001000000080006E7D2A;
defparam prom_inst_40.INIT_RAM_10 = 256'h0781FFB1FFFFFFFFC34880F1EF9C402890000001000008000007DFA700250000;
defparam prom_inst_40.INIT_RAM_11 = 256'h9FFFFFFFFC766020FFFEF318080000000000000000007EF8A02FE10FC27FBF80;
defparam prom_inst_40.INIT_RAM_12 = 256'hFF876900EB47FFE8125A00000000000000000FB780F9F664FCAFFFF801F81FFA;
defparam prom_inst_40.INIT_RAM_13 = 256'h10BBFBEEF003310000000000000000FAFA0002B006FAFFFC013F58FF28FFFDFF;
defparam prom_inst_40.INIT_RAM_14 = 256'hEFFF6D30000000000000000FF7800028000DEFFFC117F49FF2BFFFFFFFFC21E0;
defparam prom_inst_40.INIT_RAM_15 = 256'hC000000000000000F8F2800000017CFFEFCFFF39FE4BFFFFFFFF86CF82FAB8FF;
defparam prom_inst_40.INIT_RAM_16 = 256'h000000000FCF00000000044FFFA7FFF69FCF3FFFFFFFF8223E6EEE46BEFFE018;
defparam prom_inst_40.INIT_RAM_17 = 256'h003CB80000003278FFFFF7FE62F813FFFFFFFF83680E3FDCF7DEFFC67B880000;
defparam prom_inst_40.INIT_RAM_18 = 256'h000004BC8FFFFFFFE50F0C3FFFFFFFF836D0B2FF2AFDFFFCC411800000000000;
defparam prom_inst_40.INIT_RAM_19 = 256'hF1FFFFFFFE01F033FFFFFFFF03BA459FEFDF7FFFE201D480000000000003CBC0;
defparam prom_inst_40.INIT_RAM_1A = 256'hFFCD8E067FFFFFFFF03AC2282F83FFFFFE829C30000000000000FC8600000068;
defparam prom_inst_40.INIT_RAM_1B = 256'hA7FFFFFFFFC197987B827EEFFFFB630C78000000000003C4D140002F751FFFFF;
defparam prom_inst_40.INIT_RAM_1C = 256'hFFE00C99CB430EFFFFFECCB17B000000000000FE27CF200E5E23FFFFFFFDD803;
defparam prom_inst_40.INIT_RAM_1D = 256'hD7653BBEAFFFB87CEBF6000000001261F1352BBA09847FFFFFFFA980465FFFFF;
defparam prom_inst_40.INIT_RAM_1E = 256'h27D7FA0EECFAF981000040247F0D1E654020C3FFFFFFF63805C7FFFFFFFF8035;
defparam prom_inst_40.INIT_RAM_1F = 256'hFC1EF7A74300010407FC335F9D3DD07FFFFFF86280F43FFFFFFFF80329D2089E;
defparam prom_inst_40.INIT_RAM_20 = 256'h023000883BFFF0FC1F0CEE0FFFFFFF04480A47FFFFFFFFE03979B2CB4D7DFD10;
defparam prom_inst_40.INIT_RAM_21 = 256'h332FFF83204D4883FFFFFFF0CEC1047FFFFFFDFC01CD5A82AC332FF71FCDCF7F;
defparam prom_inst_40.INIT_RAM_22 = 256'h0E661A60FFFFFFFC082CF3C7FFFFFFFFF80F34A836E783FE33FD17DBF1170700;
defparam prom_inst_40.INIT_RAM_23 = 256'h1FFFFFFF81599D847FFFFFFFFF803891C07E796FD3BFB86E9FFFBFA67CFEFFFC;
defparam prom_inst_40.INIT_RAM_24 = 256'hF0185DBBC3FFFFFFFFFE03E24AD38E12FD37F18EE1FAF3BFD6FFFFFFF4180030;
defparam prom_inst_40.INIT_RAM_25 = 256'hD45FFFFFFFFFD00F8EA3EC7E8EEF3F788E7FEFFEFFFFFFFFFFF03FF807FFFFFF;
defparam prom_inst_40.INIT_RAM_26 = 256'hFFFFFD00BE230F96E09DF0E02BFCFFFFEFE7FFFFFFFFC00003FFFFFFFF8191F8;
defparam prom_inst_40.INIT_RAM_27 = 256'h01FCD6FF8F00BB0ED30FBBFFFFF7FFFFDFFFFF00023FFFFFDF4016BBBFC7FFFF;
defparam prom_inst_40.INIT_RAM_28 = 256'h7EB1F950E820B4FFFFFFFFFFFFFFFFFF800FFFFFEFF701873B085FFFFF7FFFF4;
defparam prom_inst_40.INIT_RAM_29 = 256'h06E603B3FFFFFFFFFFFFFFFFF1A7FFFFFCDB200FC1B689FFFDF6BB93C005F95A;
defparam prom_inst_40.INIT_RAM_2A = 256'h9FFFFFFFFFFFFFFFFFFFFFFE3F7C28000017F83EF3FBD0FF74000FF50DFB6348;
defparam prom_inst_40.INIT_RAM_2B = 256'hFFFFFFFFFFFDFFFFBE5100000001D100C47B6403BB80000FC9BFF7DD78E82038;
defparam prom_inst_40.INIT_RAM_2C = 256'hFFFFFD7FFCF0000000000860003E0048C08200001F22DFD199CCC001EDFFFFFF;
defparam prom_inst_40.INIT_RAM_2D = 256'hE6CC1000000000BC0000040401240A00003C97FC2C4E95000E9FFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2E = 256'h00000000000000000010000000003A47FCF6E20803F57FFFFFFFFFFFFFFFFE5E;
defparam prom_inst_40.INIT_RAM_2F = 256'h0000000000000000000001CF9FEA57E4003C8FFFFFFFFFFFFFFFFFE1EEA10000;
defparam prom_inst_40.INIT_RAM_30 = 256'h000000000001C0073A7F8600E007E67FFFFFFFFFFBF7EFE7F50C000000000000;
defparam prom_inst_40.INIT_RAM_31 = 256'h000063001D3BF9E02C00F60FFFFFFFFFFFDFFF9EDB9400000000000000000000;
defparam prom_inst_40.INIT_RAM_32 = 256'h2064E73939900360FFFFFFFFDFFC1EEF97000000000000000000000000000000;
defparam prom_inst_40.INIT_RAM_33 = 256'h482001380FFFFFFFFFE0140A0000CA00000000000000000000000000000021B3;
defparam prom_inst_40.INIT_RAM_34 = 256'hC0FFFFFFFF4C400000800000000000000000000000000000000003FFFC03B3B0;
defparam prom_inst_40.INIT_RAM_35 = 256'hF37C40000000000000000000000000000000000000000038FFF01CED08C0000F;
defparam prom_inst_40.INIT_RAM_36 = 256'h00000000000000000000000000000000000000007FFFF03AB855000B750477FF;
defparam prom_inst_40.INIT_RAM_37 = 256'h0000002000000000000000000000000003FFFF81CB4540011E013FFDD7410000;
defparam prom_inst_40.INIT_RAM_38 = 256'h2E68000000000A0020500000002BFFFC074A9BE01BD8178C1E48000000000000;
defparam prom_inst_40.INIT_RAM_39 = 256'h202252E25E7B50400000BDFFF0396E08C29F00FC000E00000000000000000020;
defparam prom_inst_40.INIT_RAM_3A = 256'hCFFFFE10000003FFFF80E6BD57FAE82F81418000000000000000007C1BDFF044;
defparam prom_inst_40.INIT_RAM_3B = 256'hC000000FFFFF833A13CB8907F80BB0000000000000000077FFFFFFAE1BFEDBDE;
defparam prom_inst_40.INIT_RAM_3C = 256'h3FFFF81E6A0B2B102A8A3600400000000000003FBB7FBFFFFECF2FE7F7FFFE80;
defparam prom_inst_40.INIT_RAM_3D = 256'h39A1655B006001000000000111680033FFFFFFF7FF9FFF7F7EFFFFFFFA10000B;
defparam prom_inst_40.INIT_RAM_3E = 256'hC04402000000000400484237BFFFFFFFFFFFFFFFFFFFFFFFFFFA000004FFFFC0;
defparam prom_inst_40.INIT_RAM_3F = 256'h00000003392E885EFF7FFFFFFFFFFFFFFFFFFFFFFFFFEE40002FFFFF00E31DF5;

pROM prom_inst_41 (
    .DO({prom_inst_41_dout_w[30:0],prom_inst_41_dout[12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_41.READ_MODE = 1'b1;
defparam prom_inst_41.BIT_WIDTH = 1;
defparam prom_inst_41.RESET_MODE = "SYNC";
defparam prom_inst_41.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFF91001FFFFFF0AC0A8BFF2A0FFFFFE57FC701FFFFFFFC000FF;
defparam prom_inst_41.INIT_RAM_01 = 256'hFFFFFFFFE8001FFFFFE4E00084FE741FFFFFE07F8301FFFFFFFC001C67FFBBFF;
defparam prom_inst_41.INIT_RAM_02 = 256'hFFC003FFFFF85840087FC8C1FFFFFE6FF8503FFFFFFFC0174F56FEEBFFFFFFFF;
defparam prom_inst_41.INIT_RAM_03 = 256'hFFFE6E400037FBE81FFFFFEEFF0700FFFFFFD000FD817FFBDFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_04 = 256'h08207EAD81FFFFFE4FF0600FFFFFF2003B3405BFF7FFFFFFFFFFFFFFFFFA011F;
defparam prom_inst_41.INIT_RAM_05 = 256'hB01FFFFFECFF0601BFFFFF8007BF80E9FF57FFFFFFFFFFFFFFFFE38FFFFFEBD2;
defparam prom_inst_41.INIT_RAM_06 = 256'hFE9FE0E01FFFFFFC00E4E027CF7D7FFFFFFFFFFFFFFFFFC3FFFFF47060041FC7;
defparam prom_inst_41.INIT_RAM_07 = 256'h03FDFFEC001ECF00FE3F177FFFFFFFFFFFFFFFFFFFFFFE45000120FD9600FFFF;
defparam prom_inst_41.INIT_RAM_08 = 256'h0003D9801F48B61FFFFFFFFFFFFFFFFFFFFFFFD13A80202FB2C037FFFFD0FE06;
defparam prom_inst_41.INIT_RAM_09 = 256'h03EF22F97FFFFFFFFFFFFFFFFFFFFFF1360701C2EA5803FFFFF84FC0200BFFF7;
defparam prom_inst_41.INIT_RAM_0A = 256'hE2FFFFFFFFFFFFFFFFFFFFFE6B96100200E9002EFFFF946806004FFC98003A24;
defparam prom_inst_41.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFC7FB84671A08B0013FFFF14B80C0017ED900070B00FDF50F;
defparam prom_inst_41.INIT_RAM_0C = 256'hFFFFFFFFF83D30C5E0288B0007BFFF34201C0037B05000F07007DF7E7F2FFFFF;
defparam prom_inst_41.INIT_RAM_0D = 256'hFE1E8B30284088B0023FFFE34001C0008200001E0700FBEFF84DFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0E = 256'h515098AE0001FFFC0000140011800001CE4C1F7DF7A50F6FFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0F = 256'h600187FE03800380003000001D6833FFFF7802C7FFFFFFFFFFFFFFFFFF91F5FA;
defparam prom_inst_41.INIT_RAM_10 = 256'hF818001800000000038A80FEFBEF0017D7FFFFFFFFFFFFFFFFF81FBF00CD0009;
defparam prom_inst_41.INIT_RAM_11 = 256'h80000000007AB001DF7DF0005F7FFFFFFFFFFFFFFFFF82F9602CA1075600407F;
defparam prom_inst_41.INIT_RAM_12 = 256'h0007B10001FFDF0003A3FFFFFFFFFFFFFFFFF0378607E86437600007FE028002;
defparam prom_inst_41.INIT_RAM_13 = 256'h1112FBC08002CEBFFFFFFFFFFFFFFF02FA0005F001F60003FEC0680038000200;
defparam prom_inst_41.INIT_RAM_14 = 256'h00002B45FFFFFFFFFFFFFFF027800020002D60003EE805800780000000003B90;
defparam prom_inst_41.INIT_RAM_15 = 256'hDFFFFFFFFFFFFFFF01F280000000540010300018005800000000073E03243F7C;
defparam prom_inst_41.INIT_RAM_16 = 256'hFFFFFFFFF017000000000AC000580007800D00000000003BB26E10FFC0000012;
defparam prom_inst_41.INIT_RAM_17 = 256'hFFC0F800000012E8000008005000F00000000003B43FFC40F80100073E77FFFF;
defparam prom_inst_41.INIT_RAM_18 = 256'h00000351800000000B000200000000003B31CFF912020000FDC67FFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_19 = 256'hD000000000F000B00000000003D2C53FE61080000FFEAB7FFFFFFFFFFFFC0FC0;
defparam prom_inst_41.INIT_RAM_1A = 256'h000B800A00000000003C9C8A3F88C80000DF708FFFFFFFFFFFFF00FE00000006;
defparam prom_inst_41.INIT_RAM_1B = 256'hE00000000001E5E2E376A310001913EF87FFFFFFFFFFFC06F3000012FB000000;
defparam prom_inst_41.INIT_RAM_1C = 256'h00000F2EF936FB800000B34F6CFFFFFFFFFFFF003DD5400BAF6000000001B803;
defparam prom_inst_41.INIT_RAM_1D = 256'h7824047A500037FF5B89FFFFFFFFED9E01CF3884F5EC000000003F8076000000;
defparam prom_inst_41.INIT_RAM_1E = 256'hF02803FEF7FC067EFFFFBFDB800E3E0EADE5C000000007980740000000000039;
defparam prom_inst_41.INIT_RAM_1F = 256'hFF7EE858BCFFFEFBF8003D9F827EB0000000007D80FC000000000003CC7E1361;
defparam prom_inst_41.INIT_RAM_20 = 256'hFDCFFF77C40000E2E1F0A60000000007D80EC000000000003E68D24DDC02002F;
defparam prom_inst_41.INIT_RAM_21 = 256'hCCD00003C4A9DB8000000000BDC1EC000000000001F1A5889FECD006FFFACE00;
defparam prom_inst_41.INIT_RAM_22 = 256'h0F87F9E0000000000D1CECC000000000000FC6C82B786A00CFFEE7E80EE8F8FF;
defparam prom_inst_41.INIT_RAM_23 = 256'h0000000001FB9E4C0000000000003F19E0AB4790087FD76E0000405983010000;
defparam prom_inst_41.INIT_RAM_24 = 256'h00173DC4C0000000000003FC6AC0A1EBC18FFC7EEC050C4029000000001FFFF0;
defparam prom_inst_41.INIT_RAM_25 = 256'h2C0000000000000FF32302917A70FFA6EEF010010000000000003FF800000000;
defparam prom_inst_41.INIT_RAM_26 = 256'h00000000BFC5CC331FF60FFBCB7F80001018000000000000000000000001F7FF;
defparam prom_inst_41.INIT_RAM_27 = 256'h01FF1A2068F8E0FF6D0FB00000080000200000000000000000001C7BC2C00000;
defparam prom_inst_41.INIT_RAM_28 = 256'h813E1F0FF7E0B9C0000000000000000000000000000001FF3ED8000000000000;
defparam prom_inst_41.INIT_RAM_29 = 256'hFF5A03F80000000000000000000000000000000FC1C98000000000000005FE64;
defparam prom_inst_41.INIT_RAM_2A = 256'h800000000000000000000000000000000018D8000000000000000FF990051D39;
defparam prom_inst_41.INIT_RAM_2B = 256'h0000000000000000000000000001AB00000000000000000FF2401629C7F7A03F;
defparam prom_inst_41.INIT_RAM_2C = 256'h000000000000000000000D6000000000000000001FC9205E543FB801F8000000;
defparam prom_inst_41.INIT_RAM_2D = 256'h00000000000000BC0000000000000000003F2D035321EA800F40000000000000;
defparam prom_inst_41.INIT_RAM_2E = 256'h00000000000000000000000000003CB806211CE803F800000000000000000000;
defparam prom_inst_41.INIT_RAM_2F = 256'h0000000000000000000001F4E03DA838003E0000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_30 = 256'h0000000000000007D3817BCF0007D40000000000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_31 = 256'h000000001E4E0FFFDD00EF000000000000000000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_32 = 256'h007930E20D980360000000000000000000000000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_33 = 256'h3020413E00000000000000000000000000000000000000000000000000000000;
defparam prom_inst_41.INIT_RAM_34 = 256'hC00000000000000000000000000000000000000000000000000000000003C4C0;
defparam prom_inst_41.INIT_RAM_35 = 256'h00000000000000000000000000000000000000000000000000001F330140020F;
defparam prom_inst_41.INIT_RAM_36 = 256'h00000000000000000000000000000000000000000000003CD020001B71000000;
defparam prom_inst_41.INIT_RAM_37 = 256'h0000002000000000000000000000000000000001F24C10009F80000000000000;
defparam prom_inst_41.INIT_RAM_38 = 256'h2E68000000000A002050000000000000078D466077F000000000000000000000;
defparam prom_inst_41.INIT_RAM_39 = 256'h202252E25E7B504000000000003E7017D6BE0000000000000000000000000020;
defparam prom_inst_41.INIT_RAM_3A = 256'hCFFFFE10000000000000F8C0AFFFD80000000000000000000000007C1BDFF044;
defparam prom_inst_41.INIT_RAM_3B = 256'hC0000000000003C36C3FFD00000000000000000000000077FFFFFFAE1BFEDBDE;
defparam prom_inst_41.INIT_RAM_3C = 256'h0000001F8DC665B000000000000000000000003FBB7FBFFFFECF2FE7F7FFFE80;
defparam prom_inst_41.INIT_RAM_3D = 256'h3E3B1E27000000000000000111680033FFFFFFF7FF9FFF7F7EFFFFFFFA100000;
defparam prom_inst_41.INIT_RAM_3E = 256'hC00000000000000400484237BFFFFFFFFFFFFFFFFFFFFFFFFFFA000000000000;
defparam prom_inst_41.INIT_RAM_3F = 256'h00000003392E885EFF7FFFFFFFFFFFFFFFFFFFFFFFFFEE400000000000FC1C37;

pROM prom_inst_42 (
    .DO({prom_inst_42_dout_w[30:0],prom_inst_42_dout[13]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_42.READ_MODE = 1'b1;
defparam prom_inst_42.BIT_WIDTH = 1;
defparam prom_inst_42.RESET_MODE = "SYNC";
defparam prom_inst_42.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFD1001FFFFFFF8405710019FFFFFFFEFFF8FFFFFFFFFFFFF18;
defparam prom_inst_42.INIT_RAM_01 = 256'hFFFFFFFFE8001FFFFFF80021C200B3FFFFFFFDFFF8FFFFFFFFFFFFE508004FFF;
defparam prom_inst_42.INIT_RAM_02 = 256'hFF4003FFFFFE22010840163FFFFFFFBFFF8FFFFFFFFFFFE820A9013FFFFFFFFF;
defparam prom_inst_42.INIT_RAM_03 = 256'hFFFFA12004100027FFFFFFF1FFF8FFFFFFFFFFFF107C8004FFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_04 = 256'h000000947FFFFFFF3FFF9FFFFFFFFFFFC30BF64007FFFFFFFFFFFFFFFFFE007F;
defparam prom_inst_42.INIT_RAM_05 = 256'h8FFFFFFFFFFFF9FFFFFFFFFFF8387F67009FFFFFFFFFFFFFFFFFF00FFFFFF800;
defparam prom_inst_42.INIT_RAM_06 = 256'hFF7FFF1FFFFFFFFFFF060FD8B4867FFFFFFFFFFFFFFFFFFFFFFFFE010000001A;
defparam prom_inst_42.INIT_RAM_07 = 256'hFFFFFFFFFFE0C0FF03D0B9FFFFFFFFFFFFFFFFFFFFFFFFC17800000631FFFFFF;
defparam prom_inst_42.INIT_RAM_08 = 256'hFFFC1C7FC03F49AFFFFFFFFFFFFFFFFFFFFFFFE13D800400463FFFFFFFEBFFF1;
defparam prom_inst_42.INIT_RAM_09 = 256'hFC00FD03BFFFFFFFFFFFFFFFFFFFFFFD37F300C00CC7FFFFFFFFBFFF5FFFFFFF;
defparam prom_inst_42.INIT_RAM_0A = 256'h24FFFFFFFFFFFFFFFFFFFFFFABE9B00A10B8FFFFFFFFF3FFF9FFFFFFFFFFC09B;
defparam prom_inst_42.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFBF47AE7F20D8FFFFFFFFEBFFF3FFFFFFFFFF8087F000270;
defparam prom_inst_42.INIT_RAM_0C = 256'hFFFFFFFFFF5FDF3DFFF8D8FFFFFFFFC3FFE3FFFFFFFFFF010FF800018333FFFF;
defparam prom_inst_42.INIT_RAM_0D = 256'hFFE0FFB7FBBF8D8FFFFFFFFC3FFEBFFFFFFFFFE038FE000007BD5FFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0E = 256'h7FAF78F9FFFFFFFFD7FFE3FFFFFFFFFE0733C000005AFE7FFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0F = 256'h1FFFFFFFFD7FFC7FFFFFFFFFE137CC000003F981FFFFFFFFFFFFFFFFFFFE0AF2;
defparam prom_inst_42.INIT_RAM_10 = 256'hFFE7FFC7FFFFFFFFFC1E7F0000007FE0EFFFFFFFFFFFFFFFFFFFF05F00BAFF8D;
defparam prom_inst_42.INIT_RAM_11 = 256'h7FFFFFFFFF834FFF00000FFF83BFFFFFFFFFFFFFFFFFFD07E02EDEF791FFFFFF;
defparam prom_inst_42.INIT_RAM_12 = 256'hFFF834FF3A0000FFFC08FFFFFFFFFFFFFFFFFFC87DFFFF9BF91FFFFFFFFC7FFD;
defparam prom_inst_42.INIT_RAM_13 = 256'hEEE4001F7FFC63BFFFFFFFFFFFFFFFFD05FFFDCFFF11FFFFFFFF87FFC7FFFFFF;
defparam prom_inst_42.INIT_RAM_14 = 256'hFFFFD8DBFFFFFFFFFFFFFFFFC87FFFDFFFFB1FFFFFFFFA7FF87FFFFFFFFFC3CF;
defparam prom_inst_42.INIT_RAM_15 = 256'h3FFFFFFFFFFFFFFFFE0D7FFFFFFFB3FFFFFFFFE7FFC7FFFFFFFFF83E7CDBC003;
defparam prom_inst_42.INIT_RAM_16 = 256'hFFFFFFFFFFE8FFFFFFFFF23FFFFFFFF87FF0FFFFFFFFFFC3B191EF803FFFFFBC;
defparam prom_inst_42.INIT_RAM_17 = 256'hFFFF07FFFFFFFD27FFFFFFFF8FFF0FFFFFFFFFFC3C0003BD07FFFFF923FFFFFF;
defparam prom_inst_42.INIT_RAM_18 = 256'hFFFFFFA47FFFFFFFF4FFF9FFFFFFFFFFC3F02006F1FFFFFF0033FFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_19 = 256'h4FFFFFFFFF4FFF0FFFFFFFFFFC1DC24019EFFFFFF8008FFFFFFFFFFFFFFFF03F;
defparam prom_inst_42.INIT_RAM_1A = 256'hFFF47FE1FFFFFFFFFFC0E215C07737FFFFA0013FFFFFFFFFFFFFFF01FFFFFF61;
defparam prom_inst_42.INIT_RAM_1B = 256'h1FFFFFFFFFFE062804845CFFFFE6FC30FFFFFFFFFFFFFFF88E7FFFEC08FFFFFF;
defparam prom_inst_42.INIT_RAM_1C = 256'hFFFFF0312080017FFFFE7FF08FFFFFFFFFFFFFFFC2317FF7011FFFFFFFFE07FC;
defparam prom_inst_42.INIT_RAM_1D = 256'h90024015FFFFCFFF843FFFFFFFFFFFFFFE088B5FC223FFFFFFFFD07F81FFFFFF;
defparam prom_inst_42.INIT_RAM_1E = 256'hD7FFFEFEF801FFFFFFFFFFFFFFF041E7B25C3FFFFFFFF847F83FFFFFFFFFFFC1;
defparam prom_inst_42.INIT_RAM_1F = 256'hFF810FFFFFFFFFFFFFFFC1207C918FFFFFFFFF847F13FFFFFFFFFFFC0F768C00;
defparam prom_inst_42.INIT_RAM_20 = 256'hFFFFFFFFFFFFFF020E1761FFFFFFFFF847F03FFFFFFFFFFFC0743038235FFFDF;
defparam prom_inst_42.INIT_RAM_21 = 256'hFFFFFFFC068EB87FFFFFFFFF043E23FFFFFFFFFFFE01C78160117FF9FFF0307F;
defparam prom_inst_42.INIT_RAM_22 = 256'hF007F81FFFFFFFFFF683003FFFFFFFFFFFF00718068615FFBFFF0813FFFFFFFF;
defparam prom_inst_42.INIT_RAM_23 = 256'hFFFFFFFFFE086123FFFFFFFFFFFFC01EE018402FF7FFE090DFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_24 = 256'hFFE802023FFFFFFFFFFFFC0074C050043C7FFE010FFFFFFFFFFFFFFFFFE0000F;
defparam prom_inst_42.INIT_RAM_25 = 256'h63FFFFFFFFFFFFF003D30000058FFFC010EFFFFFFFFFFFFFFFFFC007FFFFFFFF;
defparam prom_inst_42.INIT_RAM_26 = 256'hFFFFFFFF40064C080061FFFC040F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000;
defparam prom_inst_42.INIT_RAM_27 = 256'hFE001E2030071FFF80F1BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE004063FFFFF;
defparam prom_inst_42.INIT_RAM_28 = 256'h80E020FFF81F437FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00C207FFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_29 = 256'hFF81FC13FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF03E047FFFFFFFFFFFFFFA007F;
defparam prom_inst_42.INIT_RAM_2A = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE047FFFFFFFFFFFFFFF001FC028007;
defparam prom_inst_42.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE08FFFFFFFFFFFFFFFFF003F00C043FF85FC0;
defparam prom_inst_42.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFF11FFFFFFFFFFFFFFFFFE00FC02073FF07FE03FFFFFF;
defparam prom_inst_42.INIT_RAM_2D = 256'hFFFFFFFFFFFFFF43FFFFFFFFFFFFFFFFFFC03F00811FF07FF03FFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0F80104FF17FC07FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFE07E02C07C1FFC17FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFF81F8180301FF803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_31 = 256'hFFFFFFFFE07E080012FF10FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_32 = 256'hFF81F0540667FD8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_33 = 256'h03DFBEC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_34 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC07C0;
defparam prom_inst_42.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03F003FFDF0;
defparam prom_inst_42.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0E383FFE48AFFFFFF;
defparam prom_inst_42.INIT_RAM_37 = 256'hFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE039B0FFF603FFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_38 = 256'hD197FFFFFFFFF5FFDFAFFFFFFFFFFFFFF80E061FF807FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_39 = 256'hDFDDAD1DA184AFBFFFFFFFFFFFC07A4026C0FFFFFFFFFFFFFFFFFFFFFFFFFFDF;
defparam prom_inst_42.INIT_RAM_3A = 256'h300001EFFFFFFFFFFFFF00E053FC17FFFFFFFFFFFFFFFFFFFFFFFF83E4200FBB;
defparam prom_inst_42.INIT_RAM_3B = 256'h3FFFFFFFFFFFFC038CAFE0FFFFFFFFFFFFFFFFFFFFFFFF8800000051E4012421;
defparam prom_inst_42.INIT_RAM_3C = 256'hFFFFFFE00E119E0FFFFFFFFFFFFFFFFFFFFFFFC0448040000130D0180800017F;
defparam prom_inst_42.INIT_RAM_3D = 256'hC03F0020FFFFFFFFFFFFFFFEEE97FFCC00000008006000808100000005EFFFFF;
defparam prom_inst_42.INIT_RAM_3E = 256'h3FFFFFFFFFFFFFFBFFB7BDC84000000000000000000000000005FFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3F = 256'hFFFFFFFCC6D177A1008000000000000000000000000011BFFFFFFFFFFF001C34;

pROM prom_inst_43 (
    .DO({prom_inst_43_dout_w[30:0],prom_inst_43_dout[14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_43.READ_MODE = 1'b1;
defparam prom_inst_43.BIT_WIDTH = 1;
defparam prom_inst_43.RESET_MODE = "SYNC";
defparam prom_inst_43.INIT_RAM_00 = 256'h00000000000000011000000000088380F005800000004000000000000000001C;
defparam prom_inst_43.INIT_RAM_01 = 256'h00000000080000000000003E3E00900000000200060000000000000700000000;
defparam prom_inst_43.INIT_RAM_02 = 256'h0040000000000001F7C012000000002000000000000000006000000000000000;
defparam prom_inst_43.INIT_RAM_03 = 256'h0000200007F002600000000000000000000000001C0000000000000000000000;
defparam prom_inst_43.INIT_RAM_04 = 256'h000000CC00000000000000000000000003800400000000000000000000020000;
defparam prom_inst_43.INIT_RAM_05 = 256'h8000000000000000000000000028002001000000000000000000000000000800;
defparam prom_inst_43.INIT_RAM_06 = 256'h004000000000000000040001800C0000000000000000000000000201C0000011;
defparam prom_inst_43.INIT_RAM_07 = 256'h0000000000008000060070000000000000000000000000414400000670000000;
defparam prom_inst_43.INIT_RAM_08 = 256'h00001C0020180880000000000000000000000001304004004E00000000000000;
defparam prom_inst_43.INIT_RAM_09 = 256'h04006007000000000000000000000001371F004009C0000000010000C0000000;
defparam prom_inst_43.INIT_RAM_0A = 256'h1C00000000000000000000002BC0700610980000000008000000000000000200;
defparam prom_inst_43.INIT_RAM_0B = 256'h000000000000000007F801E78B0B800000000080000000000000001800000102;
defparam prom_inst_43.INIT_RAM_0C = 256'h0000000000BE300BE008B8000000000000000000000000050000000408C00000;
defparam prom_inst_43.INIT_RAM_0D = 256'h0001C77816008B80000000000001000000000000380100001022400000000000;
defparam prom_inst_43.INIT_RAM_0E = 256'h604008980000000000000000000000000F000000004082000000000000000000;
defparam prom_inst_43.INIT_RAM_0F = 256'h00000000020000000000000001700000000002700000000000000000000101FA;
defparam prom_inst_43.INIT_RAM_10 = 256'h0010000000000000000E00400000800F00000000000000000000003F00C0008B;
defparam prom_inst_43.INIT_RAM_11 = 256'h000000000003E001000000003C0000000000000000000000E02F000FB0000000;
defparam prom_inst_43.INIT_RAM_12 = 256'h00003C000000000000F40000000000000000000003FFFE007B00000000000001;
defparam prom_inst_43.INIT_RAM_13 = 256'h00080020000390200000000000000000000003E003B000000000000000000000;
defparam prom_inst_43.INIT_RAM_14 = 256'h00000E40000000000000000010000004001300000000000000000000000003C0;
defparam prom_inst_43.INIT_RAM_15 = 256'h0000000000000000010000000000300000000040002000000000003E00002000;
defparam prom_inst_43.INIT_RAM_16 = 256'h000000000000000000000600000000020000000000000003B000008000000011;
defparam prom_inst_43.INIT_RAM_17 = 256'h00008000000000600000000000000000000000003C0000000800000020000000;
defparam prom_inst_43.INIT_RAM_18 = 256'h0000010C00000000000004000000000003F00000040000000240000000000000;
defparam prom_inst_43.INIT_RAM_19 = 256'hC00000000080000000000000001FC00000000000080480000000000000000400;
defparam prom_inst_43.INIT_RAM_1A = 256'h00040000000000000000F20000000000000008000000000000000020000000D0;
defparam prom_inst_43.INIT_RAM_1B = 256'h8000000000000788000000000000002000000000000000000180001C18000000;
defparam prom_inst_43.INIT_RAM_1C = 256'h0000003C20040000000100000800000000000000041FC00D0300000000000000;
defparam prom_inst_43.INIT_RAM_1D = 256'hCB00801000000000000000000000000000107DE7006000000000000000000000;
defparam prom_inst_43.INIT_RAM_1E = 256'h4000000101000000000000000000601E400C0000000002000200000000000001;
defparam prom_inst_43.INIT_RAM_1F = 256'h0000000000000000000001C0000380000000000400100000000000000E060600;
defparam prom_inst_43.INIT_RAM_20 = 256'h0000000000000003F008E000000000004004000000000000007CF01000000040;
defparam prom_inst_43.INIT_RAM_21 = 256'h00000000077078000000000004002000000000000001F9804000000000000000;
defparam prom_inst_43.INIT_RAM_22 = 256'h0007F800000000000080020000000000000007F8030000000000001800000000;
defparam prom_inst_43.INIT_RAM_23 = 256'h0000000000080120000000000000001F600C804000000001C000000000000000;
defparam prom_inst_43.INIT_RAM_24 = 256'h0008001200000000000000007EC02800020000001E0000000000000000000000;
defparam prom_inst_43.INIT_RAM_25 = 256'h200000000000000003E300000840000101F00000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_26 = 256'h000000000007CC0600080000001F800000000000000000000000000000001000;
defparam prom_inst_43.INIT_RAM_27 = 256'h00001E2008000000000038000000000000000000000000000000060002000000;
defparam prom_inst_43.INIT_RAM_28 = 256'h80000000002005C0000000000000000000000000000000000240000000000000;
defparam prom_inst_43.INIT_RAM_29 = 256'h000000180000000000000000000000000000000000240000000000000000007F;
defparam prom_inst_43.INIT_RAM_2A = 256'h00000000000000000000000000000000000040000000000000000001FC000080;
defparam prom_inst_43.INIT_RAM_2B = 256'h00000000000000000000000000000000000000000000000003F0040400004000;
defparam prom_inst_43.INIT_RAM_2C = 256'h0000000000000000000001000000000000000000000FC0103000000000000000;
defparam prom_inst_43.INIT_RAM_2D = 256'h0000000000000000000000000000000000003F00418000000000000000000000;
defparam prom_inst_43.INIT_RAM_2E = 256'h000000000000000000000000000000F800000010000000000000000000000000;
defparam prom_inst_43.INIT_RAM_2F = 256'h000000000000000000000007E028000200000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_30 = 256'h00000000000000001F8180004000000000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_31 = 256'h00000000007E0800000000000000000000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_32 = 256'h0001F0D504000080000000000000000000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_34 = 256'h00000000000000000000000000000000000000000000000000000000000007C0;
defparam prom_inst_43.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000003F00000000;
defparam prom_inst_43.INIT_RAM_36 = 256'h000000000000000000000000000000000000000000000000FE80000000000000;
defparam prom_inst_43.INIT_RAM_37 = 256'h000000000000000000000000000000000000000003E300010000000000000000;
defparam prom_inst_43.INIT_RAM_38 = 256'h00000000000000000000000000000000000F2200580000000000000000000000;
defparam prom_inst_43.INIT_RAM_39 = 256'h00000000000000000000000000007FA00AC00000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_3A = 256'h0000000000000000000000F2C2FE100000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_3B = 256'h0000000000000003F243F0000000000000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_3C = 256'h000000000FF02F00000000000000000000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_3D = 256'h003F006000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_43.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000001C34;

pROM prom_inst_44 (
    .DO({prom_inst_44_dout_w[30:0],prom_inst_44_dout[15]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_44.READ_MODE = 1'b1;
defparam prom_inst_44.BIT_WIDTH = 1;
defparam prom_inst_44.RESET_MODE = "SYNC";
defparam prom_inst_44.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFEEFFFFFFFFFF73C000FF87FFFFFFF9FFFDFFFFFFFFFFFFFE3;
defparam prom_inst_44.INIT_RAM_01 = 256'hFFFFFFFFF7FFFFFFFFFFFFC001FF0FFFFFFFF9FFF9FFFFFFFFFFFFF8FFFFFFFF;
defparam prom_inst_44.INIT_RAM_02 = 256'hFFBFFFFFFFFFFFFE003FE1FFFFFFFF9FFFBFFFFFFFFFFFFF9FFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_03 = 256'hFFFFDFFFF80FFC1FFFFFFFFBFFFBFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_04 = 256'hFFFFFF03FFFFFFFFBFFFBFFFFFFFFFFFFC7FFBFFFFFFFFFFFFFFFFFFFFFDFFFF;
defparam prom_inst_44.INIT_RAM_05 = 256'h7FFFFFFFF3FFFBFFFFFFFFFFFFC7FF9FFEFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF;
defparam prom_inst_44.INIT_RAM_06 = 256'hFF3FFFBFFFFFFFFFFFF9FFF07FF3FFFFFFFFFFFFFFFFFFFFFFFFFDFE3FFFFFE0;
defparam prom_inst_44.INIT_RAM_07 = 256'hFFFFFFFFFFFF3FFE01FF0FFFFFFFFFFFFFFFFFFFFFFFFFBE83FFFFF80FFFFFFF;
defparam prom_inst_44.INIT_RAM_08 = 256'hFFFFE3FFC007F07FFFFFFFFFFFFFFFFFFFFFFFFEC03FFBFF81FFFFFFFFF7FFFB;
defparam prom_inst_44.INIT_RAM_09 = 256'hF8001F80FFFFFFFFFFFFFFFFFFFFFFFEC800FF3FF03FFFFFFFFE7FFF3FFFFFFF;
defparam prom_inst_44.INIT_RAM_0A = 256'h03FFFFFFFFFFFFFFFFFFFFFFD4000FF1EF07FFFFFFFFE7FFF7FFFFFFFFFFFD7F;
defparam prom_inst_44.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFF800001804F07FFFFFFFFE7FFF7FFFFFFFFFFFE7FF8000FC;
defparam prom_inst_44.INIT_RAM_0C = 256'hFFFFFFFFFF000000000707FFFFFFFFEFFFF7FFFFFFFFFFFAFFF00003F00FFFFF;
defparam prom_inst_44.INIT_RAM_0D = 256'hFFF000000000707FFFFFFFFEFFFE7FFFFFFFFFFFC7FE00000FC03FFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0E = 256'h80000707FFFFFFFFEFFFEFFFFFFFFFFFF0FFE000003F01FFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0F = 256'hFFFFFFFFFCFFFEFFFFFFFFFFFE8FFC000007FC0FFFFFFFFFFFFFFFFFFFFE0005;
defparam prom_inst_44.INIT_RAM_10 = 256'hFFCFFFEFFFFFFFFFFFE1FF8000007FF03FFFFFFFFFFFFFFFFFFFE000FF000070;
defparam prom_inst_44.INIT_RAM_11 = 256'hFFFFFFFFFFFC1FFE00000FFFC0FFFFFFFFFFFFFFFFFFFE001FD000000FFFFFFF;
defparam prom_inst_44.INIT_RAM_12 = 256'hFFFFC3FFFC0001FFFF03FFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFDFFFC;
defparam prom_inst_44.INIT_RAM_13 = 256'hFFF0001FFFFC0FDFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFDFFFDFFFFFFF;
defparam prom_inst_44.INIT_RAM_14 = 256'hFFFFF039FFFFFFFFFFFFFFFFE00000000000FFFFFFFFFDFFFDFFFFFFFFFFFC3F;
defparam prom_inst_44.INIT_RAM_15 = 256'h1FFFFFFFFFFFFFFFFE00000000000FFFFFFFFF9FFF9FFFFFFFFFFFC1FFFFC003;
defparam prom_inst_44.INIT_RAM_16 = 256'hFFFFFFFFFFF00000000001FFFFFFFFF9FFFBFFFFFFFFFFFC4FFFFF007FFFFFE0;
defparam prom_inst_44.INIT_RAM_17 = 256'hFFFF00000000001FFFFFFFFFBFFFBFFFFFFFFFFFC3FFFFFE07FFFFF8C1FFFFFF;
defparam prom_inst_44.INIT_RAM_18 = 256'h00000003FFFFFFFFFBFFF3FFFFFFFFFFFC0FFFFFF8FFFFFF818FFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_19 = 256'h3FFFFFFFFF3FFF7FFFFFFFFFFFE03FFFFFFFFFFFF0037FFFFFFFFFFFFFFFF800;
defparam prom_inst_44.INIT_RAM_1A = 256'hFFF3FFF7FFFFFFFFFFFF01FFFFFFFFFFFF0007FFFFFFFFFFFFFFFFC000000000;
defparam prom_inst_44.INIT_RAM_1B = 256'h7FFFFFFFFFFFF807FFF9FFFFFFF0001FFFFFFFFFFFFFFFFF0000000007FFFFFF;
defparam prom_inst_44.INIT_RAM_1C = 256'hFFFFFFC01FF807FFFFFE0001F7FFFFFFFFFFFFFFF800000000FFFFFFFFFF7FFE;
defparam prom_inst_44.INIT_RAM_1D = 256'h00FF000FFFFFE0001FFFFFFFFFFFFFFFFFE00000001FFFFFFFFFE7FFEFFFFFFF;
defparam prom_inst_44.INIT_RAM_1E = 256'h3FFFFC0000FFFFFFFFFFFFFFFFFF80000003FFFFFFFFFC3FFCFFFFFFFFFFFFFE;
defparam prom_inst_44.INIT_RAM_1F = 256'h000FFFFFFFFFFFFFFFFFFE0000007FFFFFFFFFC3FFCFFFFFFFFFFFFFF001F800;
defparam prom_inst_44.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFC00001FFFFFFFFFFC3FF9FFFFFFFFFFFFFF800FE000FFFF80;
defparam prom_inst_44.INIT_RAM_21 = 256'hFFFFFFFFF80007FFFFFFFFFFC3FF9FFFFFFFFFFFFFFE007F8003FFF80000FFFF;
defparam prom_inst_44.INIT_RAM_22 = 256'hFFF807FFFFFFFFFFF87FF1FFFFFFFFFFFFFFF807FC000FFF00000FE7FFFFFFFF;
defparam prom_inst_44.INIT_RAM_23 = 256'hFFFFFFFFFF87FE1FFFFFFFFFFFFFFFE01FF0003FE00000FE3FFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_24 = 256'hFFF0FFE1FFFFFFFFFFFFFFFF813FC001FC00000FE1FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_25 = 256'h1FFFFFFFFFFFFFFFFC0CFF0007800000FE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_26 = 256'hFFFFFFFFFFF833F8003000001FE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFE;
defparam prom_inst_44.INIT_RAM_27 = 256'hFFFFE1DFF001000001FE47FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFE1FFFFFF;
defparam prom_inst_44.INIT_RAM_28 = 256'h7FC00800001FF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_29 = 256'h0003FFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFF80;
defparam prom_inst_44.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFE03FF0040;
defparam prom_inst_44.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFC0FF80200003FFF;
defparam prom_inst_44.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFF03FE0000007FFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FF800000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07FE08000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFF81FD04001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFE07E02003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_31 = 256'hFFFFFFFFFF81F0100FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_32 = 256'hFFFE0F0883FFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83F;
defparam prom_inst_44.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFFFFFF;
defparam prom_inst_44.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007FFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00FFFEFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FF87FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF801FF13FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFF003C01EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFC01F00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3C = 256'hFFFFFFFFF00FC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3D = 256'hFFC0FF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3CB;

pROM prom_inst_45 (
    .DO({prom_inst_45_dout_w[15:0],prom_inst_45_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_52),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_45.READ_MODE = 1'b1;
defparam prom_inst_45.BIT_WIDTH = 16;
defparam prom_inst_45.RESET_MODE = "SYNC";
defparam prom_inst_45.INIT_RAM_00 = 256'hAD13AD13A513AD13A513A513A513A513A513A513A513A513A513A513A513A513;
defparam prom_inst_45.INIT_RAM_01 = 256'h94709C909C919CB19CB1A4D2A4F2A4F3A4F3A513A513A513A513A513A513AD13;
defparam prom_inst_45.INIT_RAM_02 = 256'h9CD29CB294B19C9194919471947094508C2F8C0F8C0F840F8C0F8C2F94509470;
defparam prom_inst_45.INIT_RAM_03 = 256'hAD33AD33AD33AD33AD33A533A513A513A513A513A513A513A4F3A4F39CF39CD2;
defparam prom_inst_45.INIT_RAM_04 = 256'hA513AD13AD13AD33AD13AD13AD33AD33AD13AD34AD33AD33AD33AD33AD33AD34;
defparam prom_inst_45.INIT_RAM_05 = 256'hA4D2A4F2A4F2A4F2A4F2A4F3A4F3A4F3A4F3A4F3A4F3A513A4F3A513A513A513;
defparam prom_inst_45.INIT_RAM_06 = 256'h9CD29CB29CB29CB29CD29CD29CD29CD29CD29CD29CD29CD2A4D29CD2A4D29CD2;
defparam prom_inst_45.INIT_RAM_07 = 256'h9CB29CB29CD29CB29CB29CB29CB29CB29CB29CB29CD29CD29CD29CB29CB29CD2;
defparam prom_inst_45.INIT_RAM_08 = 256'h9CB29CB29CB29CD29CB29CD29CB29CB29CB29CD29CD29CB29CB29CB29CB29CD2;
defparam prom_inst_45.INIT_RAM_09 = 256'h9CB29CB29CB29CB29CD29CB29CB29CB29CD29CD29CD29CB29CD29CD29CB29CB2;
defparam prom_inst_45.INIT_RAM_0A = 256'h9CB29CD29CD29CB29CB29CD29CD29CB29CD29CD29CD29CD29CD29CD29CB29CB2;
defparam prom_inst_45.INIT_RAM_0B = 256'h9CB29CB19CB19CB29CB19CB29CB29CB19CB29CB29CB29CB29CB19CD29CB29CB2;
defparam prom_inst_45.INIT_RAM_0C = 256'h9CD29CD29CB19CD29CB19CB29CB29CB29CB29CB29CD29CB29CB29CB29CB29CB2;
defparam prom_inst_45.INIT_RAM_0D = 256'h9CD29CF2A4F39CD29CF29CD29CD29CD29CD29CB29CB29CB29CD29CB29CB29CB2;
defparam prom_inst_45.INIT_RAM_0E = 256'h9CD29CD2A4D2A4D29CD2A4D29CD29CD29CD29CD29CD29CD29CD29CD29CF29CF2;
defparam prom_inst_45.INIT_RAM_0F = 256'h9CD2A4D2A4F39CF29CF29CD2A4F3A4F39CD2A4F39CD2A4F39CF29CD29CF29CF2;
defparam prom_inst_45.INIT_RAM_10 = 256'hA4F3A4F2A4D2A4D2A4F2A4D29CD2A4F2A4D2A4F3A4D29CD2A4D2A4F3A4F3A4D2;
defparam prom_inst_45.INIT_RAM_11 = 256'hA513A4F3A4F3A4F3A513A513A513A513A4F3A513A513A513A513A4F3A4F3A4F3;
defparam prom_inst_45.INIT_RAM_12 = 256'hAD13AD13AD13AD13A513A513A513A513AD13A513A513A513A513A513A513A513;
defparam prom_inst_45.INIT_RAM_13 = 256'h9C919C919C919CB19CB19CB19CD2A4D2A4D2A4F2A4F2A4F3A513A513A513A513;
defparam prom_inst_45.INIT_RAM_14 = 256'hA513A513A4F3A513A4F3A4F39CD29CD29CD29CB29CB19CB19CB19C919C919C91;
defparam prom_inst_45.INIT_RAM_15 = 256'hAD33AD33AD33AD33AD33AD33AD33AD33AD33AD33AD13AD34A513A513A513A513;
defparam prom_inst_45.INIT_RAM_16 = 256'hA513AD13A513AD13AD13AD13AD13AD13AD13AD13AD13AD13AD13AD33AD33AD33;
defparam prom_inst_45.INIT_RAM_17 = 256'hA4D29CD29CD29CD2A4D2A4D2A4F2A4F2A4F2A4F2A4F3A4F3A4F2A4F2A4F3A4F3;
defparam prom_inst_45.INIT_RAM_18 = 256'h9CD29CD29CB29CB19CB29CB29CB29CB29CB29CD29CB29CD29CD29CD2A4D2A4D2;
defparam prom_inst_45.INIT_RAM_19 = 256'h9CB29CB19CB19CB19CB29CB29CB29CB29CB29CB29CB29CB29CB19CB29CB19CD2;
defparam prom_inst_45.INIT_RAM_1A = 256'h9CD29CB29CB29CB29CB29CB29CB29CD29CB29CB29CB29CB29CB29CD29CB29CB2;
defparam prom_inst_45.INIT_RAM_1B = 256'h9CB29CB29CB29CD29CB29CB29CD29CB29CB29CB29CB29CB29CB29CB29CB29CB2;
defparam prom_inst_45.INIT_RAM_1C = 256'h9CD29CB19CB29CB29CD29CB29CB29CB29CB29CB29CB19CB29CD29CD29CD29CD2;
defparam prom_inst_45.INIT_RAM_1D = 256'h9CB19CB29CB29CB29CB19CB29CB19CB19CB19CB19CB29CB29CB29CB29CB29CB2;
defparam prom_inst_45.INIT_RAM_1E = 256'h9CB29CB29CB19CB29CB29CB19CB29CB29CB29CB29CB29CB29CB29CB29CB29CB1;
defparam prom_inst_45.INIT_RAM_1F = 256'h9CD29CD29CD29CB29CD29CD29CD29CB29CD29CB29CD29CD29CD29CB29CB29CB2;
defparam prom_inst_45.INIT_RAM_20 = 256'h9CD29CD29CD29CD29CD2A4D29CD29CD29CD29CD29CD29CD29CD29CD29CD2A4D2;
defparam prom_inst_45.INIT_RAM_21 = 256'h9CD29CD29CD29CD29CD29CD29CD2A4D2A4D2A4D39CD29CD2A4D29CD29CD29CD2;
defparam prom_inst_45.INIT_RAM_22 = 256'hA4F2A4F3A4F3A4F2A4F2A4F2A4D2A4D2A4F2A4F2A4F2A4F29CD2A4D29CD29CD2;
defparam prom_inst_45.INIT_RAM_23 = 256'hA513A513A513A513A4F2A4F3A4F3A513A513A513A4F3A4F3A4F3A4F3A513A4F3;
defparam prom_inst_45.INIT_RAM_24 = 256'hAD13A513AD13A513A513A513AD13AD33A513AD33A513A513A513A4F3A513A513;
defparam prom_inst_45.INIT_RAM_25 = 256'hA4D29CD29CB1A4D2A4D29CD29CB19CB1A4F2A4F2A4F2A4F2A4F2A513A4F2A513;
defparam prom_inst_45.INIT_RAM_26 = 256'hAD13AD13A533A533A533A513A513A513A4F3A4F3A4F3A4F2A4F2A4F29CD29CD2;
defparam prom_inst_45.INIT_RAM_27 = 256'hAD33AD33AD33AD33AD33AD13AD33AD34AD34AD33AD33AD33AD33AD33AD33AD34;
defparam prom_inst_45.INIT_RAM_28 = 256'hA4F2A4F2A4F2A4F3A4F3A4F3A4F3AD13A513AD13AD13AD13AD13AD13AD13AD13;
defparam prom_inst_45.INIT_RAM_29 = 256'hA4D29CB29CD29CD29CD29CD29CB29CD2A4D29CD2A4F2A4D2A4F2A4F2A4F2A4F2;
defparam prom_inst_45.INIT_RAM_2A = 256'h9CB19CB29CB19CB19CB29CB29CB29CB29CB19CB29CB29CB29CB29CB19CB19CB2;
defparam prom_inst_45.INIT_RAM_2B = 256'h9CB19CB19CB29CB29CB19CB19CB29CB19CB19CB19CB19CB19CB29CB19CB19CB2;
defparam prom_inst_45.INIT_RAM_2C = 256'h9CB29CB29CB29CB29CB29CB29CB29CB29CB29CB29CB29CB29C919CB19CB19CB1;
defparam prom_inst_45.INIT_RAM_2D = 256'h9C919CB29CB29CB19CB19CB29CB19CB29CB29CB29CB29CB29CB29CB29CB29CB2;
defparam prom_inst_45.INIT_RAM_2E = 256'h9CB19CB19CB29CB19CB19CB19CB29CB19CB29CB19CB29CB19CB29CB29CB29CB1;
defparam prom_inst_45.INIT_RAM_2F = 256'h9CB19CB29CB19CB29CB29CB19CB19CB29CB19CB29CB29CB19CB19CB29CB29CB1;
defparam prom_inst_45.INIT_RAM_30 = 256'h9CB19CB29CB19CB29CB19CB19CB19CB19CB19CB19CB19CB19C919C919CB29CB2;
defparam prom_inst_45.INIT_RAM_31 = 256'h9CD29CD29CD29CD29CB29CD29CB29CD29CD29CB29CD29CB29CB29CB29CB29CB2;
defparam prom_inst_45.INIT_RAM_32 = 256'h9CD29CD29CD29CD29CD29CD29CD29CD29CD29CD29CD29CD29CD29CD29CD29CD2;
defparam prom_inst_45.INIT_RAM_33 = 256'h9CD29CD29CD29CD29CD29CD29CD29CD29CD2A4D29CD29CD29CD29CD29CD2A4D2;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_5 (
  .Q(dff_q_5),
  .D(dff_q_4),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_6 (
  .Q(dff_q_6),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_7 (
  .Q(dff_q_7),
  .D(dff_q_6),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_8 (
  .Q(dff_q_8),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_9 (
  .Q(dff_q_9),
  .D(dff_q_8),
  .CLK(clk),
  .CE(oce)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(promx9_inst_0_dout[0]),
  .I1(promx9_inst_1_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(promx9_inst_2_dout[0]),
  .I1(promx9_inst_3_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(promx9_inst_4_dout[0]),
  .I1(promx9_inst_5_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(promx9_inst_6_dout[0]),
  .I1(promx9_inst_7_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(promx9_inst_8_dout[0]),
  .I1(promx9_inst_9_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(promx9_inst_10_dout[0]),
  .I1(promx9_inst_11_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(promx9_inst_12_dout[0]),
  .I1(promx9_inst_13_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(promx9_inst_14_dout[0]),
  .I1(promx9_inst_15_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(promx9_inst_30_dout[0]),
  .I1(promx9_inst_31_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(promx9_inst_32_dout[0]),
  .I1(promx9_inst_33_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(promx9_inst_34_dout[0]),
  .I1(promx9_inst_35_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(promx9_inst_36_dout[0]),
  .I1(promx9_inst_37_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(dff_q_7)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_27),
  .I1(mux_o_28),
  .S0(dff_q_7)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_29),
  .I1(mux_o_30),
  .S0(dff_q_7)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_31),
  .I1(mux_o_32),
  .S0(dff_q_7)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(dff_q_7)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_7)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(dff_q_5)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(dff_q_5)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_5)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_3)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_47),
  .I1(prom_inst_45_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_51 (
  .O(dout[0]),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_1)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(promx9_inst_0_dout[1]),
  .I1(promx9_inst_1_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(promx9_inst_2_dout[1]),
  .I1(promx9_inst_3_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(promx9_inst_4_dout[1]),
  .I1(promx9_inst_5_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(promx9_inst_6_dout[1]),
  .I1(promx9_inst_7_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(promx9_inst_8_dout[1]),
  .I1(promx9_inst_9_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(promx9_inst_10_dout[1]),
  .I1(promx9_inst_11_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(promx9_inst_12_dout[1]),
  .I1(promx9_inst_13_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(promx9_inst_14_dout[1]),
  .I1(promx9_inst_15_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(promx9_inst_30_dout[1]),
  .I1(promx9_inst_31_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(promx9_inst_32_dout[1]),
  .I1(promx9_inst_33_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(promx9_inst_34_dout[1]),
  .I1(promx9_inst_35_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(promx9_inst_36_dout[1]),
  .I1(promx9_inst_37_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_7)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_7)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_7)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(dff_q_7)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_7)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(dff_q_7)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_5)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(dff_q_5)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(dff_q_5)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_97),
  .I1(mux_o_98),
  .S0(dff_q_3)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_99),
  .I1(prom_inst_45_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_103 (
  .O(dout[1]),
  .I0(mux_o_101),
  .I1(mux_o_102),
  .S0(dff_q_1)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(promx9_inst_0_dout[2]),
  .I1(promx9_inst_1_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(promx9_inst_2_dout[2]),
  .I1(promx9_inst_3_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(promx9_inst_4_dout[2]),
  .I1(promx9_inst_5_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(promx9_inst_6_dout[2]),
  .I1(promx9_inst_7_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(promx9_inst_8_dout[2]),
  .I1(promx9_inst_9_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(promx9_inst_10_dout[2]),
  .I1(promx9_inst_11_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(promx9_inst_12_dout[2]),
  .I1(promx9_inst_13_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(promx9_inst_14_dout[2]),
  .I1(promx9_inst_15_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(promx9_inst_30_dout[2]),
  .I1(promx9_inst_31_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(promx9_inst_32_dout[2]),
  .I1(promx9_inst_33_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(promx9_inst_34_dout[2]),
  .I1(promx9_inst_35_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(promx9_inst_36_dout[2]),
  .I1(promx9_inst_37_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(mux_o_129),
  .I1(mux_o_130),
  .S0(dff_q_7)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_131),
  .I1(mux_o_132),
  .S0(dff_q_7)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(dff_q_7)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_7)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_7)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(dff_q_7)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(dff_q_5)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(dff_q_5)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(dff_q_5)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(mux_o_149),
  .I1(mux_o_150),
  .S0(dff_q_3)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(mux_o_151),
  .I1(prom_inst_45_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_155 (
  .O(dout[2]),
  .I0(mux_o_153),
  .I1(mux_o_154),
  .S0(dff_q_1)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(promx9_inst_0_dout[3]),
  .I1(promx9_inst_1_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(promx9_inst_2_dout[3]),
  .I1(promx9_inst_3_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(promx9_inst_4_dout[3]),
  .I1(promx9_inst_5_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(promx9_inst_6_dout[3]),
  .I1(promx9_inst_7_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(promx9_inst_8_dout[3]),
  .I1(promx9_inst_9_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(promx9_inst_10_dout[3]),
  .I1(promx9_inst_11_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(promx9_inst_12_dout[3]),
  .I1(promx9_inst_13_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(promx9_inst_14_dout[3]),
  .I1(promx9_inst_15_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(promx9_inst_30_dout[3]),
  .I1(promx9_inst_31_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(promx9_inst_32_dout[3]),
  .I1(promx9_inst_33_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(promx9_inst_34_dout[3]),
  .I1(promx9_inst_35_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(promx9_inst_36_dout[3]),
  .I1(promx9_inst_37_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_7)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(dff_q_7)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(mux_o_185),
  .I1(mux_o_186),
  .S0(dff_q_7)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(mux_o_187),
  .I1(mux_o_188),
  .S0(dff_q_7)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(dff_q_7)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(dff_q_7)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(dff_q_5)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_5)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_5)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(dff_q_3)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_203),
  .I1(prom_inst_45_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_207 (
  .O(dout[3]),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_1)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(promx9_inst_0_dout[4]),
  .I1(promx9_inst_1_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(promx9_inst_2_dout[4]),
  .I1(promx9_inst_3_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(promx9_inst_4_dout[4]),
  .I1(promx9_inst_5_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(promx9_inst_6_dout[4]),
  .I1(promx9_inst_7_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(promx9_inst_8_dout[4]),
  .I1(promx9_inst_9_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(promx9_inst_10_dout[4]),
  .I1(promx9_inst_11_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(promx9_inst_12_dout[4]),
  .I1(promx9_inst_13_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(promx9_inst_14_dout[4]),
  .I1(promx9_inst_15_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(promx9_inst_30_dout[4]),
  .I1(promx9_inst_31_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(promx9_inst_32_dout[4]),
  .I1(promx9_inst_33_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(promx9_inst_34_dout[4]),
  .I1(promx9_inst_35_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(promx9_inst_36_dout[4]),
  .I1(promx9_inst_37_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_7)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_7)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_7)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(dff_q_7)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(dff_q_7)
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(dff_q_7)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(mux_o_246),
  .I1(mux_o_247),
  .S0(dff_q_5)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(dff_q_5)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(dff_q_5)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(mux_o_253),
  .I1(mux_o_254),
  .S0(dff_q_3)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(mux_o_255),
  .I1(prom_inst_45_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_259 (
  .O(dout[4]),
  .I0(mux_o_257),
  .I1(mux_o_258),
  .S0(dff_q_1)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(promx9_inst_0_dout[5]),
  .I1(promx9_inst_1_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(promx9_inst_2_dout[5]),
  .I1(promx9_inst_3_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(promx9_inst_4_dout[5]),
  .I1(promx9_inst_5_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(promx9_inst_6_dout[5]),
  .I1(promx9_inst_7_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(promx9_inst_8_dout[5]),
  .I1(promx9_inst_9_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(promx9_inst_10_dout[5]),
  .I1(promx9_inst_11_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(promx9_inst_12_dout[5]),
  .I1(promx9_inst_13_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(promx9_inst_14_dout[5]),
  .I1(promx9_inst_15_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(promx9_inst_30_dout[5]),
  .I1(promx9_inst_31_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(promx9_inst_32_dout[5]),
  .I1(promx9_inst_33_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(promx9_inst_34_dout[5]),
  .I1(promx9_inst_35_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(promx9_inst_36_dout[5]),
  .I1(promx9_inst_37_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_285),
  .I1(mux_o_286),
  .S0(dff_q_7)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_7)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_7)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_7)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(mux_o_293),
  .I1(mux_o_294),
  .S0(dff_q_7)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_295),
  .I1(mux_o_296),
  .S0(dff_q_7)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(dff_q_5)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(dff_q_5)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(dff_q_5)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(dff_q_3)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(mux_o_307),
  .I1(prom_inst_45_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_311 (
  .O(dout[5]),
  .I0(mux_o_309),
  .I1(mux_o_310),
  .S0(dff_q_1)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(promx9_inst_0_dout[6]),
  .I1(promx9_inst_1_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(promx9_inst_2_dout[6]),
  .I1(promx9_inst_3_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(promx9_inst_4_dout[6]),
  .I1(promx9_inst_5_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(promx9_inst_6_dout[6]),
  .I1(promx9_inst_7_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(promx9_inst_8_dout[6]),
  .I1(promx9_inst_9_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(promx9_inst_10_dout[6]),
  .I1(promx9_inst_11_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(promx9_inst_12_dout[6]),
  .I1(promx9_inst_13_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(promx9_inst_14_dout[6]),
  .I1(promx9_inst_15_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(promx9_inst_30_dout[6]),
  .I1(promx9_inst_31_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(promx9_inst_32_dout[6]),
  .I1(promx9_inst_33_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(promx9_inst_34_dout[6]),
  .I1(promx9_inst_35_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(promx9_inst_36_dout[6]),
  .I1(promx9_inst_37_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(mux_o_337),
  .I1(mux_o_338),
  .S0(dff_q_7)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(mux_o_339),
  .I1(mux_o_340),
  .S0(dff_q_7)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(mux_o_341),
  .I1(mux_o_342),
  .S0(dff_q_7)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(dff_q_7)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_7)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_7)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(dff_q_5)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(dff_q_5)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(dff_q_5)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_3)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_359),
  .I1(prom_inst_45_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_363 (
  .O(dout[6]),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(dff_q_1)
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(promx9_inst_0_dout[7]),
  .I1(promx9_inst_1_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(promx9_inst_2_dout[7]),
  .I1(promx9_inst_3_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(promx9_inst_4_dout[7]),
  .I1(promx9_inst_5_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(promx9_inst_6_dout[7]),
  .I1(promx9_inst_7_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(promx9_inst_8_dout[7]),
  .I1(promx9_inst_9_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(promx9_inst_10_dout[7]),
  .I1(promx9_inst_11_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(promx9_inst_12_dout[7]),
  .I1(promx9_inst_13_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(promx9_inst_14_dout[7]),
  .I1(promx9_inst_15_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(promx9_inst_30_dout[7]),
  .I1(promx9_inst_31_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(promx9_inst_32_dout[7]),
  .I1(promx9_inst_33_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(promx9_inst_34_dout[7]),
  .I1(promx9_inst_35_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(promx9_inst_36_dout[7]),
  .I1(promx9_inst_37_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(mux_o_389),
  .I1(mux_o_390),
  .S0(dff_q_7)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(mux_o_391),
  .I1(mux_o_392),
  .S0(dff_q_7)
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(mux_o_393),
  .I1(mux_o_394),
  .S0(dff_q_7)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(mux_o_395),
  .I1(mux_o_396),
  .S0(dff_q_7)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(mux_o_397),
  .I1(mux_o_398),
  .S0(dff_q_7)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(mux_o_399),
  .I1(mux_o_400),
  .S0(dff_q_7)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(dff_q_5)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(mux_o_404),
  .I1(mux_o_405),
  .S0(dff_q_5)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(mux_o_406),
  .I1(mux_o_407),
  .S0(dff_q_5)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(dff_q_3)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_411),
  .I1(prom_inst_45_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_415 (
  .O(dout[7]),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_1)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(promx9_inst_0_dout[8]),
  .I1(promx9_inst_1_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(promx9_inst_2_dout[8]),
  .I1(promx9_inst_3_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(promx9_inst_4_dout[8]),
  .I1(promx9_inst_5_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(promx9_inst_6_dout[8]),
  .I1(promx9_inst_7_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(promx9_inst_8_dout[8]),
  .I1(promx9_inst_9_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(promx9_inst_10_dout[8]),
  .I1(promx9_inst_11_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(promx9_inst_12_dout[8]),
  .I1(promx9_inst_13_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(promx9_inst_14_dout[8]),
  .I1(promx9_inst_15_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(promx9_inst_30_dout[8]),
  .I1(promx9_inst_31_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(promx9_inst_32_dout[8]),
  .I1(promx9_inst_33_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(promx9_inst_34_dout[8]),
  .I1(promx9_inst_35_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(promx9_inst_36_dout[8]),
  .I1(promx9_inst_37_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(dff_q_7)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(dff_q_7)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(dff_q_7)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(dff_q_7)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_449),
  .I1(mux_o_450),
  .S0(dff_q_7)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_451),
  .I1(mux_o_452),
  .S0(dff_q_7)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_454),
  .I1(mux_o_455),
  .S0(dff_q_5)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(dff_q_5)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_458),
  .I1(mux_o_459),
  .S0(dff_q_5)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(mux_o_461),
  .I1(mux_o_462),
  .S0(dff_q_3)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(mux_o_463),
  .I1(prom_inst_45_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_467 (
  .O(dout[8]),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_1)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(prom_inst_16_dout[9]),
  .I1(prom_inst_17_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(prom_inst_38_dout[9]),
  .I1(prom_inst_45_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_486 (
  .O(dout[9]),
  .I0(mux_o_484),
  .I1(mux_o_485),
  .S0(dff_q_1)
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(prom_inst_18_dout[10]),
  .I1(prom_inst_19_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(prom_inst_39_dout[10]),
  .I1(prom_inst_45_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_505 (
  .O(dout[10]),
  .I0(mux_o_503),
  .I1(mux_o_504),
  .S0(dff_q_1)
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(prom_inst_20_dout[11]),
  .I1(prom_inst_21_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(prom_inst_40_dout[11]),
  .I1(prom_inst_45_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_524 (
  .O(dout[11]),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(dff_q_1)
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(prom_inst_22_dout[12]),
  .I1(prom_inst_23_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(prom_inst_41_dout[12]),
  .I1(prom_inst_45_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_543 (
  .O(dout[12]),
  .I0(mux_o_541),
  .I1(mux_o_542),
  .S0(dff_q_1)
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(prom_inst_24_dout[13]),
  .I1(prom_inst_25_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(prom_inst_42_dout[13]),
  .I1(prom_inst_45_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_562 (
  .O(dout[13]),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(dff_q_1)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(prom_inst_26_dout[14]),
  .I1(prom_inst_27_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(prom_inst_43_dout[14]),
  .I1(prom_inst_45_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_581 (
  .O(dout[14]),
  .I0(mux_o_579),
  .I1(mux_o_580),
  .S0(dff_q_1)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(prom_inst_28_dout[15]),
  .I1(prom_inst_29_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(prom_inst_44_dout[15]),
  .I1(prom_inst_45_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_600 (
  .O(dout[15]),
  .I0(mux_o_598),
  .I1(mux_o_599),
  .S0(dff_q_1)
);
endmodule //Gowin_pROM5
