//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Thu Aug 31 18:35:44 2023

module Gowin_pROM3 (dout, clk, oce, ce, reset, ad);//binary slika

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [18:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [0:0] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [0:0] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [0:0] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [0:0] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [0:0] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [0:0] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [0:0] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [0:0] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [0:0] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [0:0] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [0:0] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [0:0] prom_inst_15_dout;
wire [30:0] prom_inst_16_dout_w;
wire [0:0] prom_inst_16_dout;
wire [30:0] prom_inst_17_dout_w;
wire [0:0] prom_inst_17_dout;
wire [30:0] prom_inst_18_dout_w;
wire [0:0] prom_inst_18_dout;
wire [30:0] prom_inst_19_dout_w;
wire [0:0] prom_inst_19_dout;
wire [30:0] prom_inst_20_dout_w;
wire [0:0] prom_inst_20_dout;
wire [30:0] prom_inst_21_dout_w;
wire [0:0] prom_inst_21_dout;
wire [30:0] prom_inst_22_dout_w;
wire [0:0] prom_inst_22_dout;
wire [30:0] prom_inst_23_dout_w;
wire [0:0] prom_inst_23_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;

LUT5 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_0.INIT = 32'h00000001;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(lut_f_0)
);
defparam lut_inst_1.INIT = 4'h8;
LUT5 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_2.INIT = 32'h00000002;
LUT2 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(lut_f_2)
);
defparam lut_inst_3.INIT = 4'h8;
LUT5 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_4.INIT = 32'h00000004;
LUT2 lut_inst_5 (
  .F(lut_f_5),
  .I0(ce),
  .I1(lut_f_4)
);
defparam lut_inst_5.INIT = 4'h8;
LUT5 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_6.INIT = 32'h00000008;
LUT2 lut_inst_7 (
  .F(lut_f_7),
  .I0(ce),
  .I1(lut_f_6)
);
defparam lut_inst_7.INIT = 4'h8;
LUT5 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_8.INIT = 32'h00000010;
LUT2 lut_inst_9 (
  .F(lut_f_9),
  .I0(ce),
  .I1(lut_f_8)
);
defparam lut_inst_9.INIT = 4'h8;
LUT5 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_10.INIT = 32'h00000020;
LUT2 lut_inst_11 (
  .F(lut_f_11),
  .I0(ce),
  .I1(lut_f_10)
);
defparam lut_inst_11.INIT = 4'h8;
LUT5 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_12.INIT = 32'h00000040;
LUT2 lut_inst_13 (
  .F(lut_f_13),
  .I0(ce),
  .I1(lut_f_12)
);
defparam lut_inst_13.INIT = 4'h8;
LUT5 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_14.INIT = 32'h00000080;
LUT2 lut_inst_15 (
  .F(lut_f_15),
  .I0(ce),
  .I1(lut_f_14)
);
defparam lut_inst_15.INIT = 4'h8;
LUT5 lut_inst_16 (
  .F(lut_f_16),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_16.INIT = 32'h00000100;
LUT2 lut_inst_17 (
  .F(lut_f_17),
  .I0(ce),
  .I1(lut_f_16)
);
defparam lut_inst_17.INIT = 4'h8;
LUT5 lut_inst_18 (
  .F(lut_f_18),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_18.INIT = 32'h00000200;
LUT2 lut_inst_19 (
  .F(lut_f_19),
  .I0(ce),
  .I1(lut_f_18)
);
defparam lut_inst_19.INIT = 4'h8;
LUT5 lut_inst_20 (
  .F(lut_f_20),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_20.INIT = 32'h00000400;
LUT2 lut_inst_21 (
  .F(lut_f_21),
  .I0(ce),
  .I1(lut_f_20)
);
defparam lut_inst_21.INIT = 4'h8;
LUT5 lut_inst_22 (
  .F(lut_f_22),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_22.INIT = 32'h00000800;
LUT2 lut_inst_23 (
  .F(lut_f_23),
  .I0(ce),
  .I1(lut_f_22)
);
defparam lut_inst_23.INIT = 4'h8;
LUT5 lut_inst_24 (
  .F(lut_f_24),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_24.INIT = 32'h00001000;
LUT2 lut_inst_25 (
  .F(lut_f_25),
  .I0(ce),
  .I1(lut_f_24)
);
defparam lut_inst_25.INIT = 4'h8;
LUT5 lut_inst_26 (
  .F(lut_f_26),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_26.INIT = 32'h00002000;
LUT2 lut_inst_27 (
  .F(lut_f_27),
  .I0(ce),
  .I1(lut_f_26)
);
defparam lut_inst_27.INIT = 4'h8;
LUT5 lut_inst_28 (
  .F(lut_f_28),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_28.INIT = 32'h00004000;
LUT2 lut_inst_29 (
  .F(lut_f_29),
  .I0(ce),
  .I1(lut_f_28)
);
defparam lut_inst_29.INIT = 4'h8;
LUT5 lut_inst_30 (
  .F(lut_f_30),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_30.INIT = 32'h00008000;
LUT2 lut_inst_31 (
  .F(lut_f_31),
  .I0(ce),
  .I1(lut_f_30)
);
defparam lut_inst_31.INIT = 4'h8;
LUT5 lut_inst_32 (
  .F(lut_f_32),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_32.INIT = 32'h00010000;
LUT2 lut_inst_33 (
  .F(lut_f_33),
  .I0(ce),
  .I1(lut_f_32)
);
defparam lut_inst_33.INIT = 4'h8;
LUT5 lut_inst_34 (
  .F(lut_f_34),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_34.INIT = 32'h00020000;
LUT2 lut_inst_35 (
  .F(lut_f_35),
  .I0(ce),
  .I1(lut_f_34)
);
defparam lut_inst_35.INIT = 4'h8;
LUT5 lut_inst_36 (
  .F(lut_f_36),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_36.INIT = 32'h00040000;
LUT2 lut_inst_37 (
  .F(lut_f_37),
  .I0(ce),
  .I1(lut_f_36)
);
defparam lut_inst_37.INIT = 4'h8;
LUT5 lut_inst_38 (
  .F(lut_f_38),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_38.INIT = 32'h00080000;
LUT2 lut_inst_39 (
  .F(lut_f_39),
  .I0(ce),
  .I1(lut_f_38)
);
defparam lut_inst_39.INIT = 4'h8;
LUT5 lut_inst_40 (
  .F(lut_f_40),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_40.INIT = 32'h00100000;
LUT2 lut_inst_41 (
  .F(lut_f_41),
  .I0(ce),
  .I1(lut_f_40)
);
defparam lut_inst_41.INIT = 4'h8;
LUT5 lut_inst_42 (
  .F(lut_f_42),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_42.INIT = 32'h00200000;
LUT2 lut_inst_43 (
  .F(lut_f_43),
  .I0(ce),
  .I1(lut_f_42)
);
defparam lut_inst_43.INIT = 4'h8;
LUT5 lut_inst_44 (
  .F(lut_f_44),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_44.INIT = 32'h00400000;
LUT2 lut_inst_45 (
  .F(lut_f_45),
  .I0(ce),
  .I1(lut_f_44)
);
defparam lut_inst_45.INIT = 4'h8;
LUT5 lut_inst_46 (
  .F(lut_f_46),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_46.INIT = 32'h00800000;
LUT2 lut_inst_47 (
  .F(lut_f_47),
  .I0(ce),
  .I1(lut_f_46)
);
defparam lut_inst_47.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFF99FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_10 = 256'hFFFE3807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FC003;
defparam prom_inst_2.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0F0F81FFFFFFFF;
defparam prom_inst_2.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1A = 256'hFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007FFE0FFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1D = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC007FFF87FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF300FFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803FFFFFF;
defparam prom_inst_2.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFB281FFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003FFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_26 = 256'hFFFFFFDE0FFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_29 = 256'h7FFFFFE001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_2.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2C = 256'h0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFF00;
defparam prom_inst_2.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_30 = 256'hFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFF8000001FFFF;
defparam prom_inst_2.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_33 = 256'hFFFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000FFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_36 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE040000007FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam prom_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFF;
defparam prom_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFF80000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFC00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hFC007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_02 = 256'hF800000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFF;
defparam prom_inst_3.INIT_RAM_05 = 256'h00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFF3E00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000;
defparam prom_inst_3.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_09 = 256'hFFFFFFFFFFE3E00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFF;
defparam prom_inst_3.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0C = 256'hFF83E00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0F = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000001FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFF03E000;
defparam prom_inst_3.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFC03E0003FFFFFFF;
defparam prom_inst_3.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_16 = 256'hFFFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFF803F0007FFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_18 = 256'hFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_19 = 256'hFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFE003F001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1B = 256'hFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC003F003F9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001F;
defparam prom_inst_3.INIT_RAM_1E = 256'h0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFF0003F00FE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
defparam prom_inst_3.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000F8FFFFFFF;
defparam prom_inst_3.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_22 = 256'hFFFFFFFE0001F01FC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000001F;
defparam prom_inst_3.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FC3FFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_25 = 256'h0001F03F81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000FFFFFFFFF;
defparam prom_inst_3.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FC0FFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_3.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_28 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80007C07FFFFFFFFFFFFFFFFFFFF00001F8FE;
defparam prom_inst_3.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFC0007E00FFFFFFFFFFFFFFFFFFFE00001F9FC01FFFFFF;
defparam prom_inst_3.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFF0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFFFF8003E003FFFFFFFFFFFFFFFFFFC00001FFF001FFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_31 = 256'hFFFFFFFFFFF80000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_32 = 256'hFFFFE003E001FFFFFFFFFFFFFFFFFFC00001FFE001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_34 = 256'hFFFC0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_35 = 256'hF0003FFFFFFFFFFFFFFFFFC00001FFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003;
defparam prom_inst_3.INIT_RAM_37 = 256'h000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFC00001FF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800;
defparam prom_inst_3.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFC01F0001FFF;
defparam prom_inst_3.INIT_RAM_3A = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3B = 256'hFFFFFFC00001FE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7F01F00003FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3E = 256'h0001FC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000007FFFFFF;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1FC1F80001FFFFFFFFFFFFFF8FC0;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_9),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_01 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE07F0F80000FFFFFFFFFFFFFF0FC00003FC00;
defparam prom_inst_4.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFE01FEFC0000FFFFFFFFFFFFFC0FC0000FF80001FFFFFF;
defparam prom_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_08 = 256'hFFFFFFFFFFFF00FFFC00007FFFFFFFFFFFF80FC0001FF00001FFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0A = 256'hFFC3FFFFFFFFFFF000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0B = 256'hFFFF003FFC00007F7FFFFFFFFFF00FC0003FF00001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0D = 256'hFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0E = 256'hFE00007F1FFFFFFFFFC00FE000FFF00001FFFFFFFFFFFFFFFFFFFFFDFF00FFFF;
defparam prom_inst_4.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800F;
defparam prom_inst_4.INIT_RAM_10 = 256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_11 = 256'h07FFFFFFFF800FE001FDF00003FFFFFFFFFFFFFFFFFFFFE01E007F3FFFFFFFFE;
defparam prom_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FF00003F;
defparam prom_inst_4.INIT_RAM_13 = 256'h0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_14 = 256'hFE0007E007F0F00007FFFFFFFFFFFFFFFFFFFF800C003807FFFFFFFF00000000;
defparam prom_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FF80003F01FFFFFF;
defparam prom_inst_4.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_17 = 256'h0FE0F0000FFFFFFFFFFFFFFFFFFFFF8000000003FFFFFFFF800000000003FFFF;
defparam prom_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FC0003F807FFFFFFC0007E0;
defparam prom_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1A = 256'h1FFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFFC00000000003FFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FE0003F801FFFFFF00007E03FC0F000;
defparam prom_inst_4.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFE000000000001E3FFFFFFE00000000000FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFE0001FF8001F8007FFFFE00007E07F00F0007FFFFFFF;
defparam prom_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_20 = 256'hFFFC00000000000000FFFFFFF800000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_21 = 256'hFFFFFFFFFFFFE0001FFE001F8001FFFFC00007E1FE00F800F1FFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_23 = 256'h00000000007FFFFFF800000000005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_24 = 256'hFFFFF0000FDF801FC0007FFF000007FFF800F801E1FFFFFFFFFFFFFFFFF80000;
defparam prom_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_26 = 256'h003FFFFFFE00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_27 = 256'h0FC7E00FC0001FFE000007FFF000F807C1FFFFFFFFFFFFFFFFF8000000000000;
defparam prom_inst_4.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam prom_inst_4.INIT_RAM_29 = 256'hFF000000008047FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2A = 256'hC00007FC000003FFE000F80F01FFFFFFFFFFFFFFFFF0000000000000003FFFFF;
defparam prom_inst_4.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FC1F80F;
defparam prom_inst_4.INIT_RAM_2C = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2D = 256'h000003FF8000F81E01FFFFFFFFFFFFFFFFF000001E00000000100FFFFF800000;
defparam prom_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007C07E0FC00003FC;
defparam prom_inst_4.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_30 = 256'h0000F87C01FFFFFFFFFFFFFFFF0000003FFFC000000007FFFFC00000000001FF;
defparam prom_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007E01F87E00001FC000003FF;
defparam prom_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_33 = 256'h01FFFFFFFFFFFFFFFE000023FFFFF000000003FFFFE00000080000FFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007E00FE7E00000FE000003FC0000F8F0;
defparam prom_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFC00007FFFFFFE00000003FFFFF008000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFE003F003FFF00000FE000007F80000FBE001FFFFFF;
defparam prom_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_39 = 256'hF80000FFFFFFFFF8000003FFFFF800000000001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFF803F000FFF00000FE00000FF80000FFC001FFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01;
defparam prom_inst_4.INIT_RAM_3C = 256'hFFFFFFFC000003FFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3D = 256'hFFFFFFFE03F0007FF00000FE00001FF00000FF8001FFFFFFFFFFFFFFF80003FF;
defparam prom_inst_4.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFF;
defparam prom_inst_4.INIT_RAM_3F = 256'h000000FFFFFF000000000027FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_11),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h81F8001FF800007F00003FF00000FF0001FFFFFFFFFFFFFFF8000FFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFF0003FFFFFFFFFFFFE7F;
defparam prom_inst_5.INIT_RAM_02 = 256'hFFFF808000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_03 = 256'hFC00007F0000FFF00000FE0001FFFFFFFFFFFFFFF8001FFFFFFFFFFFF800001F;
defparam prom_inst_5.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FFFF0001FFFFFFFFFFFFE1FE1F80007;
defparam prom_inst_5.INIT_RAM_05 = 256'h10000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_06 = 256'h0001FFF80001FC0001FFFFFFFFFFFFFFF0003FFFFFFFFFFFFF000007FFFFC000;
defparam prom_inst_5.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFE000FFFF0001FFFF8FFFFFFFE07F9F80001FF00007F;
defparam prom_inst_5.INIT_RAM_08 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_09 = 256'h0003FC0001FFFFFFFFFFFFFFC0003FFFFFFFFFFFFF800007FFFFE02800000000;
defparam prom_inst_5.INIT_RAM_0A = 256'hFFFFFFFFFFFFFC0007FFF0001FFFC01FFFFFFF01FFFC0001FFC0007F0003FBF8;
defparam prom_inst_5.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0C = 256'h03FFFFFFFFFFFFFF80007FFFFFFFFFFFFFE00003FFFFF000000100003FFFFFFF;
defparam prom_inst_5.INIT_RAM_0D = 256'hFFFFFC0003FFF0001FFF800FFFFFFF00FFFC0000FFE0007F000FE3F80007FC00;
defparam prom_inst_5.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0F = 256'hFFFFFFFF8000FFFFFFFFFFFFFFF00003FFFFF804000000001FFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_10 = 256'h03FFF0001FFF0007FFFFFF801FFC0000FFF8003F801FC1F8000FFC0007FFFFFF;
defparam prom_inst_5.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_5.INIT_RAM_12 = 256'h0003FFFFFFFFFFFFFFFC0003FFFFFC00000000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_13 = 256'h1FFF0007FFFFFF8007FE0000FFFE003F807F01F8003F7C000FFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFF000;
defparam prom_inst_5.INIT_RAM_15 = 256'hFFFFFFFFFFFF0001FFFFFE000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_16 = 256'hFFFFFF8001FF00007CFF803F80FE01F8007C7C001FFFFFFFFFFFFFFF0003FFFF;
defparam prom_inst_5.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFF8001FFF0003;
defparam prom_inst_5.INIT_RAM_18 = 256'hFFFF00001FFFFF000400000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_19 = 256'h00FF80007C7FE03F81F801F800F87C003FFFFFFFFFFFFFFF0003FFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFC003FFF0003FFFFFFC0;
defparam prom_inst_5.INIT_RAM_1B = 256'h07FFFF800000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1C = 256'h7C1FF81F87F001FC03E07C00FFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFF8000;
defparam prom_inst_5.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC0FFE0003FFFF00FFFF0003FFFFFFC0007FE000;
defparam prom_inst_5.INIT_RAM_1E = 256'h00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1F = 256'hCFC001FC07C07C01FFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFF800003FFFFC0;
defparam prom_inst_5.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFF001FF0003FFFFC0FFFF0003FFFFFFE0003FF8003C07FE1F;
defparam prom_inst_5.INIT_RAM_21 = 256'h001E0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_22 = 256'h1F807C03FFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFFFFC00003FFFFE000000000;
defparam prom_inst_5.INIT_RAM_23 = 256'hFFFFFFFFE000FFC001FFFFE0FFFF0007FFFFFFE0001FFE003E01FF9FFF8001FC;
defparam prom_inst_5.INIT_RAM_24 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFF00003FFFFF00000000000000000;
defparam prom_inst_5.INIT_RAM_26 = 256'hE0007FF800FFFFE07FFF8007FFFFFFF0001FFF803E007FFFFF0000FC3E007C0F;
defparam prom_inst_5.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_28 = 256'hFFFFFFFC001FFFFFFFFFFFFFFFFFFC0003FFFFFC0000000000000000007FFFFF;
defparam prom_inst_5.INIT_RAM_29 = 256'h003FFFE03FFF801FFFFFFFF0000FFFE03E001FFFFC0000FC7C007C1FFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFF;
defparam prom_inst_5.INIT_RAM_2B = 256'h001FFFFFFFFFFFFFFFFFFF0003FFFFFE0000000000000000000FFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2C = 256'h1FFFC0FFFFFFFFF8000F8FF83F0007FFF80000FFF8007C3FFFFFFFFFFFFFFFFC;
defparam prom_inst_5.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFF801FFFE0;
defparam prom_inst_5.INIT_RAM_2E = 256'hFFFFFFFFFFFFFF0003FFFFFF00000000000000000001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2F = 256'hFFFFFFFE000FC3FE1F0001FFE00000FFE0007CFFFFFFFFFFFFFFFFFC000FFFFF;
defparam prom_inst_5.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFC007FFE00FFF81FF;
defparam prom_inst_5.INIT_RAM_31 = 256'hFFFFFF8003FFFFFF800000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_32 = 256'h8007C0FF1F00007FC00000FFC0003FFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFC001FFE007FD01FFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_34 = 256'h01FFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_35 = 256'hFF00003FC00000FF80003FFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFF80;
defparam prom_inst_5.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE00001FFE0007FC001F001FFFFFFFFFFE007C07F;
defparam prom_inst_5.INIT_RAM_37 = 256'hE000000000002000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_38 = 256'hC00000FF00003FFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFC000FFFFFF;
defparam prom_inst_5.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFF000007FF0000000000001FFFFFFFFFFF007E01FFF80001F;
defparam prom_inst_5.INIT_RAM_3A = 256'h00008000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3B = 256'h00003FFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFC0007FFFFFF0000000;
defparam prom_inst_5.INIT_RAM_3C = 256'hFFFFFFFFF800001FF0000000000003FFFFFFFFFFFC03E007FF80000FC00000FE;
defparam prom_inst_5.INIT_RAM_3D = 256'h0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFE000FFFFFFFFFFFFFFFFFFFC0007FFFFFF800000000140000;
defparam prom_inst_5.INIT_RAM_3F = 256'hFF000003F8000000000003FFFFFFFFFFFF03E001FF80000FC00001FE00007FFF;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_13),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_01 = 256'hFFFFFFFF0007FFFFFFFFFFFFFFFFFFC0007FFFFFFC000000006000000000003F;
defparam prom_inst_6.INIT_RAM_02 = 256'h00000000000003FFFFFFFFFFFFC1F0007FC0000FC00003FE00007FFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000;
defparam prom_inst_6.INIT_RAM_04 = 256'h0007FFFFFFFFFFFFFFFFFFC0007FFFFFFE000000020000000000000FFFFFFFFF;
defparam prom_inst_6.INIT_RAM_05 = 256'h000003FFFFFFFFFFFFF1F0001FE0000FE0000FFE0000FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
defparam prom_inst_6.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFE000FFFFFFFF0000000400000000000007FFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_08 = 256'hFFFFFFFFFFFDF00007F00007E0001FFE0003FFFFFFFFFFFFFFFFFFFF0003FFFF;
defparam prom_inst_6.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000003FF;
defparam prom_inst_6.INIT_RAM_0A = 256'hFFFFFFE000FFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0B = 256'hFFFFF80003FC0007E0007F3E0007FFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000007FFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0D = 256'h01FFFFFFFFC000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0E = 256'h03FF0007E000FC3F000FFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_6.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000007FFFFFFFFFFFFFFF800;
defparam prom_inst_6.INIT_RAM_10 = 256'hFFE080000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_11 = 256'hF003F83F003FFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFE001FFFFFF;
defparam prom_inst_6.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFC0000000000000007FFFFFFFFFFFFFFF80003FFC007;
defparam prom_inst_6.INIT_RAM_13 = 256'h00000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_14 = 256'h007FFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFC000FFFFFFFFF00000;
defparam prom_inst_6.INIT_RAM_15 = 256'hFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFFC0001FFF007F007F01F;
defparam prom_inst_6.INIT_RAM_16 = 256'h000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFC000FFFFFFFFF8000000000000;
defparam prom_inst_6.INIT_RAM_18 = 256'hFFFFFF8000000000000007FFFFFFFFFFFFFFFF0001F3F803F00FC01F00FFFFFF;
defparam prom_inst_6.INIT_RAM_19 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1A = 256'hFFFFFFFFC0003FFFFFFFFFFFFFFFFFC000FFFFFFFFF800000000000000000000;
defparam prom_inst_6.INIT_RAM_1B = 256'h00000000000009FFFFFFFFFFFFFFFFC001F8FE03F03F801F01FFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_6.INIT_RAM_1D = 256'hE0003FFFFFFFFFFFFFFFFF8000FFFFFFFFFC000000000000000000000FFFFFFF;
defparam prom_inst_6.INIT_RAM_1E = 256'h00000E7FFFFFFFFFFFFFFFF001F83F83F07F001F07FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000;
defparam prom_inst_6.INIT_RAM_20 = 256'hFFFFFFFFFFFFFE0001FFFFFFFFFE000000000000000000000FFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFC00F80FE3F8FC001F0FFFFFFFFFFFFFFFFFFFFFFFF0003FFF;
defparam prom_inst_6.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000003FF;
defparam prom_inst_6.INIT_RAM_23 = 256'hFFFFF80001FFFFFFFFFF0000000000000000000007FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_24 = 256'hFFFFFFFE00F803F3FFF8001F1FFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_26 = 256'h03FFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_27 = 256'h80FC00FFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFF000;
defparam prom_inst_6.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803C00000000003FFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_29 = 256'hFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_2A = 256'hFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFF0000FFFFFFF;
defparam prom_inst_6.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFE07C003F;
defparam prom_inst_6.INIT_RAM_2C = 256'h000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFE0003FFFFFFFFFFF0000;
defparam prom_inst_6.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFF800000000000FFFFFFFFFFFFFFFFFF87C000FFF80000F;
defparam prom_inst_6.INIT_RAM_2F = 256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFE0003FFFFFFFFFFF000000000000;
defparam prom_inst_6.INIT_RAM_31 = 256'hFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFE7E0003FF00000FFFFFFFFF;
defparam prom_inst_6.INIT_RAM_32 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_33 = 256'hFFFFFFFFFE0000FFFFFFFFFFFFFFC0003FFFFFFFFFFF00000000000000000000;
defparam prom_inst_6.INIT_RAM_34 = 256'hFFE0000000000003FFFFFFFFFFFFFFFFFFFE0000FE00000FFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_36 = 256'hFF0000FFFFFFFFFFFFFF00007FFFFFFFFFFE0000000000000000000000FFFFFF;
defparam prom_inst_6.INIT_RAM_37 = 256'h00000001FFFFFFFFFFFFFFFFFFFE00007E00001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam prom_inst_6.INIT_RAM_39 = 256'hFFFFFFFFFFFE00007FFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFE00003E00003FFFFFFFFFFFFFFFFFFFFFFFFFFF8000FF;
defparam prom_inst_6.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001;
defparam prom_inst_6.INIT_RAM_3C = 256'hFFFC0000FFFFFFFFFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3D = 256'hFFFFFFFFFFFF00003F00007FFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000FFFFFFFF;
defparam prom_inst_6.INIT_RAM_3F = 256'hFFFFFFFFFFFC0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_15),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'hFFFF80003F0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFF80003;
defparam prom_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_02 = 256'hFFFE0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_03 = 256'h1F0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFC00000FFFFFFFFF;
defparam prom_inst_7.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000007FFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_7.INIT_RAM_05 = 256'h000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFF000001FFFFFFFFFFFFE0000;
defparam prom_inst_7.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFF800000000000003FFFFFFFFFFFFFFFFFFFF0001F0007FF;
defparam prom_inst_7.INIT_RAM_08 = 256'h00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFE000001FFFFFFFFFFFFE000000000000;
defparam prom_inst_7.INIT_RAM_0A = 256'hFFFFFFFFFF000000000000001FFFFFFFFFFFFFFFFFFFFC001F800FFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0B = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFFF00007FFFFFFFFC000003FFFFFFFFFFFFF00000000000000000000;
defparam prom_inst_7.INIT_RAM_0D = 256'hFF000000000000001FFFFFFFFFFFFFFFFFFFFF001F803FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0F = 256'hFFFC0007FFFFFFF0C000007FFFFFFFFFFFFF0000000000000000000000FFFFFF;
defparam prom_inst_7.INIT_RAM_10 = 256'h000000000FFFFFFFFFFFFFFFFFFFFFC01F807FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
defparam prom_inst_7.INIT_RAM_12 = 256'hFFFFFFC0000000FFFFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_13 = 256'h0FFFFFFFFFFFFFFFFFFFFFF00F80FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003;
defparam prom_inst_7.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000;
defparam prom_inst_7.INIT_RAM_15 = 256'h000001FFFFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFC0F83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003C7FFFF00;
defparam prom_inst_7.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000FFFFFFF;
defparam prom_inst_7.INIT_RAM_18 = 256'hFFFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_19 = 256'hFFFFFFFF0FC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000FE0E0000001FFF;
defparam prom_inst_7.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1B = 256'hFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1C = 256'hCFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007800000001FFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1E = 256'h000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000002000000003FFFFFFFFFFFFFFFFE000;
defparam prom_inst_7.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_21 = 256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFFFF00000000000;
defparam prom_inst_7.INIT_RAM_23 = 256'hFFFFFFFFFF800000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_24 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_25 = 256'hFFFFFFFFFFFF800000000000003FFFFFFFFFFFFFFFFFF0000000000000000000;
defparam prom_inst_7.INIT_RAM_26 = 256'hFFC00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_28 = 256'hFFFFE0000000000007FFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFF;
defparam prom_inst_7.INIT_RAM_29 = 256'h000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam prom_inst_7.INIT_RAM_2B = 256'h000001801FFFFFFFFFFFFFFFFFFFFE00000000000000000001FFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC20;
defparam prom_inst_7.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000;
defparam prom_inst_7.INIT_RAM_2E = 256'h3FFFFFFFFFFFFFFFFFFFFE00000000000000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000C0;
defparam prom_inst_7.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000001FFFFFFFF;
defparam prom_inst_7.INIT_RAM_31 = 256'hFFFFFFFFFFFFFF00000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001E0FFFFFFFF;
defparam prom_inst_7.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000001FFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_34 = 256'hFFFFFF80000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000009FFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_37 = 256'h000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00C013FFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_7.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3A = 256'h0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFF87F81FFFFFFFFFFFFFFFFFFFFFFFFFE000000000;
defparam prom_inst_7.INIT_RAM_3C = 256'hFFFFFFFFFFFC00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3D = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000;
defparam prom_inst_7.INIT_RAM_3F = 256'hFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_17),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b0;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000003FFFFFF;
defparam prom_inst_8.INIT_RAM_02 = 256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000;
defparam prom_inst_8.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000F93;
defparam prom_inst_8.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF000000000000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000007F87FFFFFFFF;
defparam prom_inst_8.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFF800000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000001FFFCFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0D = 256'hFFFFFFFFE00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFDFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_10 = 256'hF800000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFDC7FFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_13 = 256'h00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000;
defparam prom_inst_8.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFDFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_16 = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000;
defparam prom_inst_8.INIT_RAM_18 = 256'hFFFFFFF9FFFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000005FFFFF;
defparam prom_inst_8.INIT_RAM_1B = 256'h3FFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_8.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800F;
defparam prom_inst_8.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFF;
defparam prom_inst_8.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFF80200000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF820003FFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFF0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01800FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_29 = 256'hFFFFFFF8000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF00403FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2C = 256'h080000000006FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_8.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2F = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
defparam prom_inst_8.INIT_RAM_31 = 256'hFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFF;
defparam prom_inst_8.INIT_RAM_34 = 256'hFE00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000003FFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF87FFFF;
defparam prom_inst_8.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFC008000000005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_19),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b0;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_02 = 256'hFFFFFFFFFE010000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01FFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_05 = 256'hFF808000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_08 = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE00300FFFFFFFFFFFFFFFFFFFFFFFFFC02000;
defparam prom_inst_9.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFE0300000C0005F;
defparam prom_inst_9.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_0F = 256'hFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFF010000100001FFFFFFFFF;
defparam prom_inst_9.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_12 = 256'hFFE00000FFFFFFFFFFFFFFFFFFFFFFFFFFF808000000000FFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC060004000007FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE60007F;
defparam prom_inst_9.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFE040000000005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0781FFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01FFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1B = 256'hFFFFFFFFFFFF030000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE27FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1E = 256'hFFFF8080000080107FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_21 = 256'h000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFF9C7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0C0;
defparam prom_inst_9.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFE1E000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_24 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_25 = 256'hFFFFFFFFFFFF10FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE06000000000;
defparam prom_inst_9.INIT_RAM_26 = 256'hFFFFFFFFFFFE3E0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_28 = 256'hFF0C1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF028010000003FFFFFFF;
defparam prom_inst_9.INIT_RAM_29 = 256'hFFFE3C0E01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8080000000007FFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2C = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE307FFFF;
defparam prom_inst_9.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE781F;
defparam prom_inst_9.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC083000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2F = 256'hFFFFFFFFFFF800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC081FFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F83E01FFFFFF;
defparam prom_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFE060000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_32 = 256'hFF000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1F07C01FFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFFFFFF028008000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_35 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFE00807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1E07C03FFFFFFFFFFFFFFFC000000;
defparam prom_inst_9.INIT_RAM_37 = 256'hFFFFFF8180000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC3C0F803FFFFFFFFFFFFFFF800000003FFFFFF;
defparam prom_inst_9.INIT_RAM_3A = 256'h40000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_3B = 256'hFFFFFFC107FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_9.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFE7C1F001FFFFFFFFFFFFFFF0000000007FFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_3D = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000;
defparam prom_inst_9.INIT_RAM_3F = 256'hFFFFFFFFFFCF83E003FFFFFFFFFFFFFFE0000000001FFFFFFFFFFFFFFFFFFC03;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_21),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b0;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF020400000000FFFFF;
defparam prom_inst_10.INIT_RAM_02 = 256'hFF0F07C007FFFFFFFFFFFFFFC00000000007FFFFFFFFFFFFFFFF847FFFFFFFFF;
defparam prom_inst_10.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8180000000007FFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_05 = 256'h1FFFFFFFFFFFFFFFC00000000003FFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1F0F80;
defparam prom_inst_10.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0E0000000003FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_08 = 256'hFFFFFFFF800000000001FFFFFFFFFFFFFFC67FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3E1F803FFFFFFF;
defparam prom_inst_10.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFE000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0B = 256'h800000000000FFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3C3F003FFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFF020020000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0E = 256'h00007FFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC787E003FFFFFFFFFFFFFFF80000000;
defparam prom_inst_10.INIT_RAM_10 = 256'hFFFFFFFF8100000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_11 = 256'hFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80FFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC7878007FFFFFFFFFFFFFFF0000000000007FFF;
defparam prom_inst_10.INIT_RAM_13 = 256'hC1C0002000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_14 = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFC00F020FFFFFFFFFFFFFFFF0000000000007FFFFFFFFFF0;
defparam prom_inst_10.INIT_RAM_16 = 256'h00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFE0600000;
defparam prom_inst_10.INIT_RAM_18 = 256'hFFFFFFFFF801F003FFFFFFFFFFFFFFFF0000000000007FFFFFFFFFC1FFFFFFFF;
defparam prom_inst_10.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1A = 256'hFFFFFFF800000007FFE0000000000FFFFFFFFFFFFFFFFFFFF028020000001FFF;
defparam prom_inst_10.INIT_RAM_1B = 256'hF8004003FFFFFFFFFFFFFFFF0000000000007FFFFFFFFC0FFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1D = 256'h000000000000000000007FFFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFF000000000000FFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFF000;
defparam prom_inst_10.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000003;
defparam prom_inst_10.INIT_RAM_20 = 256'h0007FFF001FFFFFFFFFFFFFFFFFFFFFFFC100000000003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_21 = 256'hFFFFFFFF000000000000FFFFFFFF83FFFFFFFFFFFFFFFFFFFFE00003FFFFFC00;
defparam prom_inst_10.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FFFFFFFF;
defparam prom_inst_10.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE080000000001FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_24 = 256'h000000000000FFFFFFFE1FFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFF020000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_27 = 256'h0001FFFFFFF07FFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1E0003FFFFFFFFFFFFFFFFF80000000;
defparam prom_inst_10.INIT_RAM_29 = 256'hFFFFFFFFFF8300000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_2A = 256'hFFC3FFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFF803C00FFFFFFFFFFFFFFFFFF800000000003FFFF;
defparam prom_inst_10.INIT_RAM_2C = 256'hFFC1A0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_2D = 256'hFFFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFF000E01FFFFFFFFFFFFFFFFFF800000000003FFFFFE0FFFFF;
defparam prom_inst_10.INIT_RAM_2F = 256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_30 = 256'hFFFFC01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0C000;
defparam prom_inst_10.INIT_RAM_31 = 256'hFFFFFFFF000007FFFFFFFFFFFFFFFFFFC00000000007FFFFF87FFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF020000000000F;
defparam prom_inst_10.INIT_RAM_34 = 256'h00000FFFFFFFFFFFFFFFFFFFC0000000000FFFFFE1FFFFFFFFFFFFFFFFFE01FF;
defparam prom_inst_10.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_10.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFF;
defparam prom_inst_10.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFE0000000001FFFFF87FFFFFFFFFFFFFFFFF80FFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00001FFF;
defparam prom_inst_10.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC080000000001FFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_3A = 256'hFFFFFFFFE0000000007FFFFC1FFFFFFFFFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_3D = 256'hF000000000FFFFF8FFFFFFFFFFFFFFFFFE03FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_23),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b0;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'h01FFFFE3FFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFF0000000;
defparam prom_inst_11.INIT_RAM_02 = 256'hFFFFFFFFFFFFC000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFFFFFFFF800000003FFFF9F;
defparam prom_inst_11.INIT_RAM_05 = 256'hFFFFE000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_06 = 256'hFFFFFFFE03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFF80000000FFFFE3FFFFFFFFF;
defparam prom_inst_11.INIT_RAM_08 = 256'h000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_09 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_11.INIT_RAM_0A = 256'hFFFFFF800007FFFFFFFFFFFFFFFFFFFFFC0000001FFFF8FFFFFFFFFFFFFFFFF8;
defparam prom_inst_11.INIT_RAM_0B = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000;
defparam prom_inst_11.INIT_RAM_0D = 256'h000FFFFFFFFFFFFFFFFFFFFFFC0000007FFFE1FFFFFFFFFFFFFFFFC07FFFFFFF;
defparam prom_inst_11.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_11.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000003FFFFFF;
defparam prom_inst_11.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFE000000FFFFC7FFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FFFFF;
defparam prom_inst_11.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000001FFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_13 = 256'hFFFFFFFFFF000003FFFF1FFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_16 = 256'hFF00000FFFFC3FFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_19 = 256'hFFF8FFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFFFFF80003F;
defparam prom_inst_11.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFC000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1C = 256'hFFFFFFFFFFF80FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFC000FFFFE3FFFF;
defparam prom_inst_11.INIT_RAM_1E = 256'hFFFFFFE000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1F = 256'hFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_20 = 256'hFFFFFFFFFFFFE00000FFFFFFFFFFFFFFFFFFFFFFFFE003FFFFC7FFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_21 = 256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_11.INIT_RAM_23 = 256'hFFFFC00001FFFFFFFFFFFFFFFFFFFFFFFFF01FFFFF1FFFFFFFFFFFFFFF81FFFF;
defparam prom_inst_11.INIT_RAM_24 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000;
defparam prom_inst_11.INIT_RAM_26 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFC0FFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_11.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFF;
defparam prom_inst_11.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800003FFFFFF;
defparam prom_inst_11.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFF80FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000008000007FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_2F = 256'hFFFFFFFFF7FFFFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_32 = 256'hE7FFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_35 = 256'hFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFF;
defparam prom_inst_11.INIT_RAM_37 = 256'hFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_39 = 256'hFFFFFFFFFFF800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFF81;
defparam prom_inst_11.INIT_RAM_3A = 256'hF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3C = 256'hFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFE07FFFFFFFF;
defparam prom_inst_11.INIT_RAM_3D = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000;
defparam prom_inst_11.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFF81FFFFFFFFFFFFFFFFF;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_25),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b0;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000;
defparam prom_inst_12.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000002000001FF;
defparam prom_inst_12.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFF;
defparam prom_inst_12.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFF9FFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_08 = 256'hFFFFFFF3FFFFFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0B = 256'hFFFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;
defparam prom_inst_12.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFC000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0E = 256'hFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_10 = 256'hFFFFFFFFFFE0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_12 = 256'hFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFF0FFFF;
defparam prom_inst_12.INIT_RAM_13 = 256'hFFF0000004000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_15 = 256'hF800001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFE1FFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_16 = 256'h02000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000;
defparam prom_inst_12.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000001F;
defparam prom_inst_12.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000;
defparam prom_inst_12.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000203FFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000007FFFFFFF;
defparam prom_inst_12.INIT_RAM_1E = 256'hFFFFFFFFFFFFFC7FFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000003FFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_21 = 256'hFFFFFCFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_24 = 256'hFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF800000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF;
defparam prom_inst_12.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFC000001000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_27 = 256'hF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFF000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_29 = 256'hFFFFFFFFFFFFE0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2B = 256'hFFFFFFFE000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFE1FFFFFF;
defparam prom_inst_12.INIT_RAM_2C = 256'hFFFFF0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2E = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFE3FFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2F = 256'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_12.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800;
defparam prom_inst_12.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_32 = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FF;
defparam prom_inst_12.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000;
defparam prom_inst_12.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000FFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000003FFFFF;
defparam prom_inst_12.INIT_RAM_37 = 256'hFFFFFFFFFFFF3FFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000001FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000001FFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3A = 256'hFFFE7FFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000101FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001000000FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3D = 256'hFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFC000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFF;
defparam prom_inst_12.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_27),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b0;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_01 = 256'hFFFFFFFFFFFFFF8000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFF8;
defparam prom_inst_13.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFE0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_04 = 256'hFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFF8FFFFFFFF;
defparam prom_inst_13.INIT_RAM_05 = 256'hFFFFFFF8000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFF1FFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_08 = 256'h0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam prom_inst_13.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_13.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0B = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000001FFFF;
defparam prom_inst_13.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000;
defparam prom_inst_13.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000003FFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000004000001FFF;
defparam prom_inst_13.INIT_RAM_10 = 256'hFFFFFFFFFF8FFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000FFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_13 = 256'hFF9FFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_16 = 256'hFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFE000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFF;
defparam prom_inst_13.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1A = 256'hFFFFFFFFFFFFC000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFE3F;
defparam prom_inst_13.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFF0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1D = 256'hFFFF8000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFC3FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1E = 256'hFFFFFFFFF8000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_20 = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFC7FFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_21 = 256'hFC0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_13.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_24 = 256'h4000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFF;
defparam prom_inst_13.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000;
defparam prom_inst_13.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFF9FFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000F;
defparam prom_inst_13.INIT_RAM_29 = 256'hFFFFFFFFF3FFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000007FFFFFFFF;
defparam prom_inst_13.INIT_RAM_2C = 256'hE3FFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000003FFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2F = 256'hFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFF80000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFF;
defparam prom_inst_13.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_33 = 256'hFFFFFFFFFF00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFF8FFF;
defparam prom_inst_13.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFF0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_36 = 256'hFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFF0FFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_37 = 256'hFFFFFFFFFFF80000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_39 = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFF1FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_3A = 256'hFFFC0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000;
defparam prom_inst_13.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_3D = 256'h000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000FFFFFFF;
defparam prom_inst_13.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000;
defparam prom_inst_13.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFF3FFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_29),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b0;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000001FFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000;
defparam prom_inst_14.INIT_RAM_02 = 256'hFFFFFFFE7FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000003FFFFFF;
defparam prom_inst_14.INIT_RAM_05 = 256'hFFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE000001F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_14.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000001FFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_08 = 256'hFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFC000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0C = 256'hFFFFFFFF8000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFF1FFFF;
defparam prom_inst_14.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFF80000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0F = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFE3FFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_10 = 256'hFFFFFFFFFFFFFC0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_13 = 256'hFFFFFE0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000FF;
defparam prom_inst_14.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_16 = 256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000001FFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_14.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFE3FFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_19 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000;
defparam prom_inst_14.INIT_RAM_1B = 256'hFFFFFFE7FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001FFFF;
defparam prom_inst_14.INIT_RAM_1E = 256'hFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFC00000007FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFC7;
defparam prom_inst_14.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000FFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_21 = 256'hFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_22 = 256'hFFFFFFFFFFFFF00000000FFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000007FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_25 = 256'hFFFFC00000001FFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFE3FFFFF;
defparam prom_inst_14.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFF80000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_28 = 256'h00001FFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFE3FFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_14.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_2B = 256'hFFFE3FFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_2C = 256'hFFFFFFFE0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFF;
defparam prom_inst_14.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_2F = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000001FFFFFFE3FFF;
defparam prom_inst_14.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_31 = 256'hFFFFFFFFFFFFFF3FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_32 = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFF1FFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000;
defparam prom_inst_14.INIT_RAM_34 = 256'hFFFFFE3FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000FFFFFFF1FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001FF;
defparam prom_inst_14.INIT_RAM_37 = 256'hFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFF0000000000FFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFE7F;
defparam prom_inst_14.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000FFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_3A = 256'hF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_3B = 256'hFFFFFFFFFFE0000000000FFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFF;
defparam prom_inst_14.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_3E = 256'hFFE0000000000FFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFE3FFFFFF;
defparam prom_inst_14.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF80000000000003FFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_31),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b0;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_01 = 256'h00000FFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFE3FFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFC0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam prom_inst_15.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_04 = 256'hFFFE0FFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_05 = 256'hFFFFFFFFFE0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000FFF;
defparam prom_inst_15.INIT_RAM_06 = 256'hFFFFFFFFFFE03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_08 = 256'hFF0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000FFFFFFE0FFF;
defparam prom_inst_15.INIT_RAM_09 = 256'hFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0A = 256'hFFFFFFFFFFFFF9FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0B = 256'h0800000FFFFFFFFFFFFFFFFFFFFFFF83FFC0000000000FFFFFFC0FFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000;
defparam prom_inst_15.INIT_RAM_0D = 256'hFFFFF1FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF01FFFF;
defparam prom_inst_15.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFF01FFC0000000001FFFFFFC0FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000F;
defparam prom_inst_15.INIT_RAM_10 = 256'hFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_11 = 256'hFFFFFFFFFFFFFE00FFC0000000001FFFFFF81FFFFFFFFFFFFFFFFFFFFFFFF3FF;
defparam prom_inst_15.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFF;
defparam prom_inst_15.INIT_RAM_13 = 256'h8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_14 = 256'hFFFFFFA07FC0000000003FFFFFF81FFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_17 = 256'h7FC0000000003FFFFFF03FFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFF1FFFFFFF;
defparam prom_inst_15.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_15.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1A = 256'h00007FFFFFE03FFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFF1FFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFC000000000007FFFFFFFFFFFFFFFFFFFFFFC8FFE00000;
defparam prom_inst_15.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1D = 256'hFFE07FFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1E = 256'hFFFFFFFFFFFE000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFE000000000FFFF;
defparam prom_inst_15.INIT_RAM_1F = 256'hFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_21 = 256'hFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFC07FFF;
defparam prom_inst_15.INIT_RAM_22 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_23 = 256'hFFFFFFFFFFFFC7FFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_15.INIT_RAM_24 = 256'h0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF800000003FFFFFF80FFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_15.INIT_RAM_26 = 256'hFFFFC7FFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFF;
defparam prom_inst_15.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000FFFFFFE01FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000F;
defparam prom_inst_15.INIT_RAM_29 = 256'hFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFE0000001FFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFFCFFF;
defparam prom_inst_15.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2C = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2D = 256'hFFFFEFFFFFFF8000007FFFFFF803FFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFE;
defparam prom_inst_15.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_30 = 256'hFFFFE00003FFFFFFC007FFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFE3FFFFFFF;
defparam prom_inst_15.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFFCFFF;
defparam prom_inst_15.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_33 = 256'h1FFFFFFF800FFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFE3FFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFF000000007FFFFFFFFFFFFFFFFFFFFF0FFFFFFFFC00;
defparam prom_inst_15.INIT_RAM_35 = 256'hFFFFFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_36 = 256'h801FFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_37 = 256'hFFFFFFFFFFFFFF80000000FFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_38 = 256'hFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3A = 256'hFFFFFFE0000001FFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFE003FFFFF;
defparam prom_inst_15.INIT_RAM_3B = 256'hFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3C = 256'hFFFFFFFFFFFF9FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F;
defparam prom_inst_15.INIT_RAM_3D = 256'h000007FFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFC007FFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3E = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_15.INIT_RAM_3F = 256'hFFFF1FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFC;

pROM prom_inst_16 (
    .DO({prom_inst_16_dout_w[30:0],prom_inst_16_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_16.READ_MODE = 1'b0;
defparam prom_inst_16.BIT_WIDTH = 1;
defparam prom_inst_16.RESET_MODE = "SYNC";
defparam prom_inst_16.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_01 = 256'hFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8E001FFF;
defparam prom_inst_16.INIT_RAM_02 = 256'hFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFF81FFFFFFF;
defparam prom_inst_16.INIT_RAM_03 = 256'hFFFFFFFFFFF81FFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFF1FFF;
defparam prom_inst_16.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_05 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFF007FFFFFFFC7FFFFF;
defparam prom_inst_16.INIT_RAM_06 = 256'hFFF807FFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFC;
defparam prom_inst_16.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFF001FFFFFFFE1FFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_09 = 256'hFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFC7FFFFFFF;
defparam prom_inst_16.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC007FF;
defparam prom_inst_16.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFE0007FFFFFFE07FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0C = 256'hFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFC7FFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0E = 256'hFFFFFFFFFFFFE3FFFFFFFFC0001FFFFFFF01FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0F = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFC00;
defparam prom_inst_16.INIT_RAM_11 = 256'hFFFFC7FFFFFFFF800007FFFFFF007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFF9FFFFFFFC007FFFFFFF;
defparam prom_inst_16.INIT_RAM_14 = 256'hFFFFFF000001FFFFFF001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_15 = 256'hFFFFFFFFFFFCFFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFF;
defparam prom_inst_16.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFE7FFFFFFF801FFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_17 = 256'h00007FFFFF800FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_18 = 256'hFFFCFFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFF00;
defparam prom_inst_16.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFE00007FFFFFFCFFFFFFFF003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1A = 256'hFF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1B = 256'hFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFE0000003FFF;
defparam prom_inst_16.INIT_RAM_1C = 256'hFFFFFFFF800007FFFFFF8FFFFFFFF007FFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFF;
defparam prom_inst_16.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE3FFFFFFFFC00000007FFFFC000FF;
defparam prom_inst_16.INIT_RAM_1F = 256'h8000063FFFFF8FFFFDFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFF9;
defparam prom_inst_16.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA;
defparam prom_inst_16.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFDC7FFFFFFFF800000003FFFFC0003FFFFFFFFF;
defparam prom_inst_16.INIT_RAM_22 = 256'hFFFF87FFF9FFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFF1FFFFFFFF;
defparam prom_inst_16.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000FF;
defparam prom_inst_16.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFDC7FFFFFFFF000000000FFFFC00007FFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_25 = 256'hF3FFF01FFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFF1FFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000007FFFFF83FF;
defparam prom_inst_16.INIT_RAM_27 = 256'hFFFFFFFFFFB8FFFFFFFFE0000000003FFFE00001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF00000003FFFFF80FFE3FFF03F;
defparam prom_inst_16.INIT_RAM_2A = 256'hFF78FFFFFFFFE0000000000FFFF800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8FFFF800000000FFFFFC01FE3FFF03FFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2D = 256'hFFFFC00000000003FFFE00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2E = 256'hFFFFFFFFFFF1FFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF71FFFF;
defparam prom_inst_16.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFF1FFFF8000000007FFFF0001F1FFF03FFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_30 = 256'h00000000FFFF800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_31 = 256'hFFF3FFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF1FFFFFFFF8000;
defparam prom_inst_16.INIT_RAM_32 = 256'hFFFFFFFFF0FFFE0000000181FFFC000070FFF03FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_33 = 256'h3FFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_34 = 256'hFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000;
defparam prom_inst_16.INIT_RAM_35 = 256'hE07FFC00600000307FF8000000FFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFF;
defparam prom_inst_16.INIT_RAM_36 = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDC1FFFFFFFF0000000000000FFFF800;
defparam prom_inst_16.INIT_RAM_38 = 256'hE000000C03F80000007FF03FFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFE3;
defparam prom_inst_16.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FF000;
defparam prom_inst_16.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF807FFFFFFE00000000000003FFFE000007FFFF;
defparam prom_inst_16.INIT_RAM_3B = 256'h81B8000000FFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFC7FFFFFFFF;
defparam prom_inst_16.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00FA001E0000001;
defparam prom_inst_16.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFB807FFFFFFC00000000000000FFFF800003FFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3E = 256'h00FFE03FFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFC7FFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC007000FE000000030300000;

pROM prom_inst_17 (
    .DO({prom_inst_17_dout_w[30:0],prom_inst_17_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_35),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_17.READ_MODE = 1'b0;
defparam prom_inst_17.BIT_WIDTH = 1;
defparam prom_inst_17.RESET_MODE = "SYNC";
defparam prom_inst_17.INIT_RAM_00 = 256'hFFFFFFFFF700FFFFFFF8000000000000007FFFF00003FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FE000000006000000007FF03F;
defparam prom_inst_17.INIT_RAM_03 = 256'hF700FFFFFFF8000000000000001FFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8000007FE000000001C0000000FFF03FFFFFFFFF;
defparam prom_inst_17.INIT_RAM_06 = 256'hFFF00000000000000007FFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_07 = 256'hFFFFFFFFFFE7FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE01FFFF;
defparam prom_inst_17.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFF000000FFE00000000030000001FFF03FFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_09 = 256'h000000000007FFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0A = 256'hFFE7FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE01FFFFFFE00000;
defparam prom_inst_17.INIT_RAM_0B = 256'hFFFFFFFF000002FFE00000000000000000FFF03FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0C = 256'h0007FFFFE00407FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0D = 256'hFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCC03FFFFFFC0000000000000;
defparam prom_inst_17.INIT_RAM_0E = 256'h000005FFC00000000000000000FFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFF;
defparam prom_inst_17.INIT_RAM_0F = 256'hEC0601FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDC03FFFFFFC0000000000000000FFFFF;
defparam prom_inst_17.INIT_RAM_11 = 256'hC000000000000000007FE03FFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFF8F;
defparam prom_inst_17.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000067F;
defparam prom_inst_17.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF9807FFFFFF80000000000000001FFFFFFE0BC07F;
defparam prom_inst_17.INIT_RAM_14 = 256'h00000000007FF03FFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFF1FFFFFFFFF;
defparam prom_inst_17.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000FF00000000;
defparam prom_inst_17.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFB807FFFFFF00000000000000003FFFFFFF82F01FFFFFFFFF;
defparam prom_inst_17.INIT_RAM_17 = 256'h007FE03FFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFF1FFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000006F0000000000000000;
defparam prom_inst_17.INIT_RAM_19 = 256'hFFFFFFFFB00FFFFFFF00000000000000003FFFFFFFF03C0FFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000001E0000000000000000007FC03F;
defparam prom_inst_17.INIT_RAM_1C = 256'h300FFFFFFFE0000000000000007FFFFFFFFC1F03FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFCFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFE0000000400000000C2000000003FE03FFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1F = 256'hFFFC00000000000000FFFFFFFFFF0780FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_20 = 256'hFFFFFFFFFFCFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF701FFFFF;
defparam prom_inst_17.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFE0000000000000000FFF00000001FC07FFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_22 = 256'h0000000001FFFFFFFFFFC1E03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_23 = 256'hFF8FFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF601FFFFFFFFF0000;
defparam prom_inst_17.INIT_RAM_24 = 256'hFFFFFFFE00000000000000007FF00000000FC07FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_25 = 256'h01FFFFFFFFFFF0300FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_26 = 256'hFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF603FFFFFFFFFE00000000000;
defparam prom_inst_17.INIT_RAM_27 = 256'h00000000000000003FF000000007C07FFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFF;
defparam prom_inst_17.INIT_RAM_28 = 256'hFFFFFC0E03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_17.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF607FFFFFFFFFF8000000000003FFFFFF;
defparam prom_inst_17.INIT_RAM_2A = 256'h000000001FF000000003807FFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFC7F;
defparam prom_inst_17.INIT_RAM_2B = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000;
defparam prom_inst_17.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE07FFFFFFFFFFE000000000007FFFFFFFFFFFF01;
defparam prom_inst_17.INIT_RAM_2D = 256'h03E000000001807FFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFC7FFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000;
defparam prom_inst_17.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFC00000000007FFFFFFFFFFFFC0403FFFFF;
defparam prom_inst_17.INIT_RAM_30 = 256'h0000007FFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFF87FFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000C00000;
defparam prom_inst_17.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFF0000000000FFFFFFFFFFFFFF8001FFFE7FFFFFFFF;
defparam prom_inst_17.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000FF;
defparam prom_inst_17.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFE000000001FFFFFFFFFFFFFFE0007FFC1FFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFF1FFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000FFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_38 = 256'hFFFFFFFF800000001FFFFFFFFFFFFFFFC001FFC1FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_39 = 256'hFFFFFFFFFF3FFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFF000000000000000000000000000000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3B = 256'hE00000003FFFFFFFFFFFFFFFF0007F81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3C = 256'hFF3FFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3D = 256'hFFFFFFFF800000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3E = 256'h7FFFFFFFFFFFFFFFFE000801FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3F = 256'hFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000;

pROM prom_inst_18 (
    .DO({prom_inst_18_dout_w[30:0],prom_inst_18_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_37),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_18.READ_MODE = 1'b0;
defparam prom_inst_18.BIT_WIDTH = 1;
defparam prom_inst_18.RESET_MODE = "SYNC";
defparam prom_inst_18.INIT_RAM_00 = 256'h800000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFF;
defparam prom_inst_18.INIT_RAM_01 = 256'hFFFFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFE0000007FFFFFFF;
defparam prom_inst_18.INIT_RAM_03 = 256'h0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFE1FF;
defparam prom_inst_18.INIT_RAM_04 = 256'hF1FC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000;
defparam prom_inst_18.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_06 = 256'h00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFE3FFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000;
defparam prom_inst_18.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFF03F8003;
defparam prom_inst_18.INIT_RAM_09 = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFE3FFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000;
defparam prom_inst_18.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFE007E001FFFFFFFF;
defparam prom_inst_18.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000003FF;
defparam prom_inst_18.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFE0007C00FFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFCFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000001C0007FFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_11 = 256'hFFFFFFFFFFFFE007FFFFFFFFFFFFFFFFE0001F803FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_12 = 256'hFFFFFFFFFCFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFF800000000000000000000001E0007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_14 = 256'hFFFFF80FFFFFFFFFFFFFFFFFE00003F01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_15 = 256'hFCFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_16 = 256'hFFFFFFFFFC00000000000000000000000F000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFC000007E0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_18 = 256'hFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0F;
defparam prom_inst_18.INIT_RAM_19 = 256'hFE000000000000000000000307001FFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFF;
defparam prom_inst_18.INIT_RAM_1A = 256'hFFFFFFFFC000000FE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1C = 256'h000000000000000302001FFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFF0FFF;
defparam prom_inst_18.INIT_RAM_1D = 256'hC0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
defparam prom_inst_18.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1F = 256'h0000000388003FFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFF1FFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_20 = 256'h3FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000;
defparam prom_inst_18.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000;
defparam prom_inst_18.INIT_RAM_22 = 256'hC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFF1FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000C000000000000001;
defparam prom_inst_18.INIT_RAM_24 = 256'hFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000007FFFFFF;
defparam prom_inst_18.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000780000000000003CC0007FFF;
defparam prom_inst_18.INIT_RAM_27 = 256'hFFF8BBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000007FFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFF1FFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000310000000000006C0000FFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2A = 256'hFFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2B = 256'hFFFFFFFFF3FFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9087F;
defparam prom_inst_18.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFF000073470000000006E80001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2D = 256'hFE00FFFFFFFFFFFFFFFFFFFE00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2E = 256'hE3FFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC081FFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2F = 256'hFFFFFFFFFFFFC00027CE780000003E600003FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFE00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_31 = 256'hFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFE0003FFF;
defparam prom_inst_18.INIT_RAM_32 = 256'hFFFFF0000FDFE003804787000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFF;
defparam prom_inst_18.INIT_RAM_33 = 256'hFFFFFFFC00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFE00000FFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_35 = 256'h019DC04380EFC400000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFF87FFF;
defparam prom_inst_18.INIT_RAM_36 = 256'h00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800;
defparam prom_inst_18.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0037FFFFFF0000001FFFFFFFFFFFFFFFFFC;
defparam prom_inst_18.INIT_RAM_38 = 256'hF0E18000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF01FFFFFFFFF8FFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_39 = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003981FB;
defparam prom_inst_18.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFC0007FFFFF800000007FFFFFFFFFFFFFFFFC00000000;
defparam prom_inst_18.INIT_RAM_3B = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFE00FFFFFFFFF8FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000003B70E20000;
defparam prom_inst_18.INIT_RAM_3D = 256'hFFFFFFFFFFFFE020CFFFFFE00000001FFFFFFFFFFFFFFFF800000000001FFFFF;
defparam prom_inst_18.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFE00FFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000007760C0000000FFFFFF;

pROM prom_inst_19 (
    .DO({prom_inst_19_dout_w[30:0],prom_inst_19_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_39),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_19.READ_MODE = 1'b0;
defparam prom_inst_19.BIT_WIDTH = 1;
defparam prom_inst_19.RESET_MODE = "SYNC";
defparam prom_inst_19.INIT_RAM_00 = 256'hFFFFF01D07FFFFF000000007FFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFE00FFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_03 = 256'h81FFFFF800000001FFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_04 = 256'hFFFFFFFC01FFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC11;
defparam prom_inst_19.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_06 = 256'h000000007FFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_07 = 256'h01FFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0200FFFFFE;
defparam prom_inst_19.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFF0000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_19.INIT_RAM_09 = 256'h1FFFFFFFFFFFFFC0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0A = 256'hFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8200FFFFFF80000000;
defparam prom_inst_19.INIT_RAM_0B = 256'hFFFFFFFFFE000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01FFFFFF;
defparam prom_inst_19.INIT_RAM_0C = 256'hFFFFFFC0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC8001FFFFFC000000000FFFFFF;
defparam prom_inst_19.INIT_RAM_0E = 256'hFFC0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03FFFFFFFFC7FFFF;
defparam prom_inst_19.INIT_RAM_0F = 256'h000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC034FFFFFF0000000003FFFFFFFFFFF80;
defparam prom_inst_19.INIT_RAM_11 = 256'h0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03FFFFFFFF87FFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_12 = 256'h0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000;
defparam prom_inst_19.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE0087FFFFFC000000000FFFFFFFFFFF0000000000;
defparam prom_inst_19.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803FFFFFFFF8FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000003F;
defparam prom_inst_19.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFF8703FFFFFF0000000003FFFFFFFFFF00000000000007FFFF;
defparam prom_inst_19.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFF807FFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000003FFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_19 = 256'hFFFFFFFFE003FFFFFFC000000000FFFFFFFFFE00000000000007FFFF9FFFFFFF;
defparam prom_inst_19.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFF807FFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1C = 256'hFC01FFFFFFF0000000003FFFFFFFFC00000000000003FFFF87FFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1D = 256'hFFFFFFF007FFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1F = 256'hFFF8000000000FFFFFFFF800000000000003FFFFF3FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_20 = 256'h0FFFFFFFF80FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83FFFF;
defparam prom_inst_19.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_19.INIT_RAM_22 = 256'h000007FFFFFFF800000000000003FFFFE9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_23 = 256'hF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFE0000;
defparam prom_inst_19.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFF;
defparam prom_inst_19.INIT_RAM_25 = 256'hFFFFF000000000000003FFFFCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFF8000000001FF;
defparam prom_inst_19.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00FFFFFFFF00FFFFF;
defparam prom_inst_19.INIT_RAM_28 = 256'h000000000003FFFFCE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0F7FFFFFE0000000007FFFFFE000;
defparam prom_inst_19.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01FFFFFFFF00FFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2B = 256'h0003FFFFCF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7DFFFFFF8000000003FFFFFC00000000000;
defparam prom_inst_19.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01FFFFFFFF01FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2E = 256'hCF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFF1F3FFFFFE000000000FFFFF8000000000000003FFFF;
defparam prom_inst_19.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFC01FFFFFFFF01FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_32 = 256'hFFFFFFFFFFFFF8F9FFFFFF0000000007FFFF0000000000000003FFFFCFEFFFFF;
defparam prom_inst_19.INIT_RAM_33 = 256'hFFFFFFFFFFFFFF803FFFFFFFE01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_35 = 256'hFFFFFC3F3FFFFF8000000001FFFE0000000000000007FFFFCFF7FFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_36 = 256'hFFFFFF803FFFFFFFE01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_38 = 256'h8FFFFFE000000000FFFC0000000000000007FFFFCFFBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_39 = 256'h3FFFFFFFE01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1F;
defparam prom_inst_19.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam prom_inst_19.INIT_RAM_3B = 256'h000000007FF8000000000000000FFFFFCFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3C = 256'hE03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07E3FFFFF8;
defparam prom_inst_19.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF007FFFFFFF;
defparam prom_inst_19.INIT_RAM_3E = 256'h1FF0000000000000000FFFFFCFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FCFFFFFC00000000;

pROM prom_inst_20 (
    .DO({prom_inst_20_dout_w[30:0],prom_inst_20_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_41),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_20.READ_MODE = 1'b0;
defparam prom_inst_20.BIT_WIDTH = 1;
defparam prom_inst_20.RESET_MODE = "SYNC";
defparam prom_inst_20.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF807FFFFFFFC03FFFFF;
defparam prom_inst_20.INIT_RAM_01 = 256'h00000000000FFFFFDFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FF3FFFFF800000000FE00000;
defparam prom_inst_20.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFC03FFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_04 = 256'h000FFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFC0000000780000000000000;
defparam prom_inst_20.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_07 = 256'hC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFF0000000380000000000000001FFFFF;
defparam prom_inst_20.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFDFFFFFFC0000001C0000000000000001FFFFFC1FFFFFF;
defparam prom_inst_20.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFF0000000E0000000000000003FFFFFF07FFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_11 = 256'hFFFC3FFFFFFC00000070000000000000003FFFFFFC0FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_12 = 256'hFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_14 = 256'hFFFE00000038000000000000007FFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_15 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3007FF;
defparam prom_inst_20.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_17 = 256'h0018000000000000007FFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC03FFFFFF8000;
defparam prom_inst_20.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFF;
defparam prom_inst_20.INIT_RAM_1A = 256'h0000000000FFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80FFFFFFE000000C0000;
defparam prom_inst_20.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1D = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FFFFFF8000006000000000000;
defparam prom_inst_20.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FFFFFFE00000300000000000001FFFFFF;
defparam prom_inst_20.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFE07FFFFFF00000380000000000001FFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_27 = 256'hFFFFFFFFFFFFFF81FFFFFFC00000C0000000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2A = 256'hFFFFFFE07FFFFFF0000060000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2D = 256'h3FFFFFFC000030000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_20.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_30 = 256'h00001800000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFFFF;
defparam prom_inst_20.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_33 = 256'h000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFFC0001C00;
defparam prom_inst_20.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_36 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFFFF0000E0000000000;
defparam prom_inst_20.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFF8000700000000003FFFFFFF;
defparam prom_inst_20.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC1FFFFFFE000380000000007FFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_21 (
    .DO({prom_inst_21_dout_w[30:0],prom_inst_21_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_43),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_21.READ_MODE = 1'b0;
defparam prom_inst_21.BIT_WIDTH = 1;
defparam prom_inst_21.RESET_MODE = "SYNC";
defparam prom_inst_21.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFF07FFFFFF80018000000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_03 = 256'hFFFFFFFFFFE1FFFFFFC000C000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_06 = 256'hFFF07FFFFFF0006000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_09 = 256'hFFF0003000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FFF;
defparam prom_inst_21.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0C = 256'h00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07FFFF000018;
defparam prom_inst_21.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFF80000C0000001F;
defparam prom_inst_21.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_12 = 256'hCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFC000060000007FFFFFFFFF;
defparam prom_inst_21.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFF00006000001FFFFFFFFFF87FFFFFF;
defparam prom_inst_21.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFF1FFFF00003000007FFFFFFFFFF87FFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFE7FFE0060180001FFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1F = 256'hFFFFFFF1FFEE0781C000FFFFFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_22 = 256'h7FEE1FF0E00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_21.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_25 = 256'hE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFF;
defparam prom_inst_21.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_38 = 256'hFFFFFFFFFF8083FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3B = 256'hFFF0807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3E = 256'hFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF86017;

pROM prom_inst_22 (
    .DO({prom_inst_22_dout_w[30:0],prom_inst_22_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_45),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_22.READ_MODE = 1'b0;
defparam prom_inst_22.BIT_WIDTH = 1;
defparam prom_inst_22.RESET_MODE = "SYNC";
defparam prom_inst_22.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_01 = 256'hFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFF;
defparam prom_inst_22.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF82203FFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0080FFFFFFFFF1EFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80403FFFFFFFC3F7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFC0F8CFFFFFFF07FBFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_11 = 256'hFFFFFFFFFFFFFF8830FFFFFFC0FFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_14 = 256'hFFFFFFC9907FFFFF83FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_17 = 256'h020BFFFE4FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD;
defparam prom_inst_22.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1A = 256'h3FFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0004FFFC;
defparam prom_inst_22.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80427FFE1FFFF9FF;
defparam prom_inst_22.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8431FFF83FFFDFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFE0FFFCFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFB007FFF83FFE7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFE003FFFF07FE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2D = 256'hFFFFFFFFFFFE03FFFFC1FCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_30 = 256'hFFFF87FFFFF03BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_33 = 256'hFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFF;
defparam prom_inst_22.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_23 (
    .DO({prom_inst_23_dout_w[30:0],prom_inst_23_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_47),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_23.READ_MODE = 1'b0;
defparam prom_inst_23.BIT_WIDTH = 1;
defparam prom_inst_23.RESET_MODE = "SYNC";
defparam prom_inst_23.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[18]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[17]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(prom_inst_4_dout[0]),
  .I1(prom_inst_5_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(prom_inst_6_dout[0]),
  .I1(prom_inst_7_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(prom_inst_8_dout[0]),
  .I1(prom_inst_9_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(prom_inst_10_dout[0]),
  .I1(prom_inst_11_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(prom_inst_12_dout[0]),
  .I1(prom_inst_13_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(prom_inst_14_dout[0]),
  .I1(prom_inst_15_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(prom_inst_16_dout[0]),
  .I1(prom_inst_17_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(prom_inst_18_dout[0]),
  .I1(prom_inst_19_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(prom_inst_20_dout[0]),
  .I1(prom_inst_21_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(prom_inst_22_dout[0]),
  .I1(prom_inst_23_dout[0]),
  .S0(dff_q_4)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_3)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_3)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_3)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_3)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_2)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_2)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_2)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_1)
);
MUX2 mux_inst_23 (
  .O(dout[0]),
  .I0(mux_o_21),
  .I1(mux_o_20),
  .S0(dff_q_0)
);
endmodule //Gowin_pROM3
