//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Sat Aug 05 21:07:41 2023

module Gowin_pROM (dout, clk, oce, ce, reset, ad);//binary etf

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [18:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [0:0] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [0:0] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [0:0] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [0:0] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [0:0] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [0:0] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [0:0] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [0:0] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [0:0] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [0:0] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [0:0] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [0:0] prom_inst_15_dout;
wire [30:0] prom_inst_16_dout_w;
wire [0:0] prom_inst_16_dout;
wire [30:0] prom_inst_17_dout_w;
wire [0:0] prom_inst_17_dout;
wire [30:0] prom_inst_18_dout_w;
wire [0:0] prom_inst_18_dout;
wire [30:0] prom_inst_19_dout_w;
wire [0:0] prom_inst_19_dout;
wire [30:0] prom_inst_20_dout_w;
wire [0:0] prom_inst_20_dout;
wire [30:0] prom_inst_21_dout_w;
wire [0:0] prom_inst_21_dout;
wire [30:0] prom_inst_22_dout_w;
wire [0:0] prom_inst_22_dout;
wire [30:0] prom_inst_23_dout_w;
wire [0:0] prom_inst_23_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire dff_q_7;
wire dff_q_8;
wire dff_q_9;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;

LUT5 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_0.INIT = 32'h00000001;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(lut_f_0)
);
defparam lut_inst_1.INIT = 4'h8;
LUT5 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_2.INIT = 32'h00000002;
LUT2 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(lut_f_2)
);
defparam lut_inst_3.INIT = 4'h8;
LUT5 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_4.INIT = 32'h00000004;
LUT2 lut_inst_5 (
  .F(lut_f_5),
  .I0(ce),
  .I1(lut_f_4)
);
defparam lut_inst_5.INIT = 4'h8;
LUT5 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_6.INIT = 32'h00000008;
LUT2 lut_inst_7 (
  .F(lut_f_7),
  .I0(ce),
  .I1(lut_f_6)
);
defparam lut_inst_7.INIT = 4'h8;
LUT5 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_8.INIT = 32'h00000010;
LUT2 lut_inst_9 (
  .F(lut_f_9),
  .I0(ce),
  .I1(lut_f_8)
);
defparam lut_inst_9.INIT = 4'h8;
LUT5 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_10.INIT = 32'h00000020;
LUT2 lut_inst_11 (
  .F(lut_f_11),
  .I0(ce),
  .I1(lut_f_10)
);
defparam lut_inst_11.INIT = 4'h8;
LUT5 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_12.INIT = 32'h00000040;
LUT2 lut_inst_13 (
  .F(lut_f_13),
  .I0(ce),
  .I1(lut_f_12)
);
defparam lut_inst_13.INIT = 4'h8;
LUT5 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_14.INIT = 32'h00000080;
LUT2 lut_inst_15 (
  .F(lut_f_15),
  .I0(ce),
  .I1(lut_f_14)
);
defparam lut_inst_15.INIT = 4'h8;
LUT5 lut_inst_16 (
  .F(lut_f_16),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_16.INIT = 32'h00000100;
LUT2 lut_inst_17 (
  .F(lut_f_17),
  .I0(ce),
  .I1(lut_f_16)
);
defparam lut_inst_17.INIT = 4'h8;
LUT5 lut_inst_18 (
  .F(lut_f_18),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_18.INIT = 32'h00000200;
LUT2 lut_inst_19 (
  .F(lut_f_19),
  .I0(ce),
  .I1(lut_f_18)
);
defparam lut_inst_19.INIT = 4'h8;
LUT5 lut_inst_20 (
  .F(lut_f_20),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_20.INIT = 32'h00000400;
LUT2 lut_inst_21 (
  .F(lut_f_21),
  .I0(ce),
  .I1(lut_f_20)
);
defparam lut_inst_21.INIT = 4'h8;
LUT5 lut_inst_22 (
  .F(lut_f_22),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_22.INIT = 32'h00000800;
LUT2 lut_inst_23 (
  .F(lut_f_23),
  .I0(ce),
  .I1(lut_f_22)
);
defparam lut_inst_23.INIT = 4'h8;
LUT5 lut_inst_24 (
  .F(lut_f_24),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_24.INIT = 32'h00001000;
LUT2 lut_inst_25 (
  .F(lut_f_25),
  .I0(ce),
  .I1(lut_f_24)
);
defparam lut_inst_25.INIT = 4'h8;
LUT5 lut_inst_26 (
  .F(lut_f_26),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_26.INIT = 32'h00002000;
LUT2 lut_inst_27 (
  .F(lut_f_27),
  .I0(ce),
  .I1(lut_f_26)
);
defparam lut_inst_27.INIT = 4'h8;
LUT5 lut_inst_28 (
  .F(lut_f_28),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_28.INIT = 32'h00004000;
LUT2 lut_inst_29 (
  .F(lut_f_29),
  .I0(ce),
  .I1(lut_f_28)
);
defparam lut_inst_29.INIT = 4'h8;
LUT5 lut_inst_30 (
  .F(lut_f_30),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_30.INIT = 32'h00008000;
LUT2 lut_inst_31 (
  .F(lut_f_31),
  .I0(ce),
  .I1(lut_f_30)
);
defparam lut_inst_31.INIT = 4'h8;
LUT5 lut_inst_32 (
  .F(lut_f_32),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_32.INIT = 32'h00010000;
LUT2 lut_inst_33 (
  .F(lut_f_33),
  .I0(ce),
  .I1(lut_f_32)
);
defparam lut_inst_33.INIT = 4'h8;
LUT5 lut_inst_34 (
  .F(lut_f_34),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_34.INIT = 32'h00020000;
LUT2 lut_inst_35 (
  .F(lut_f_35),
  .I0(ce),
  .I1(lut_f_34)
);
defparam lut_inst_35.INIT = 4'h8;
LUT5 lut_inst_36 (
  .F(lut_f_36),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_36.INIT = 32'h00040000;
LUT2 lut_inst_37 (
  .F(lut_f_37),
  .I0(ce),
  .I1(lut_f_36)
);
defparam lut_inst_37.INIT = 4'h8;
LUT5 lut_inst_38 (
  .F(lut_f_38),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_38.INIT = 32'h00080000;
LUT2 lut_inst_39 (
  .F(lut_f_39),
  .I0(ce),
  .I1(lut_f_38)
);
defparam lut_inst_39.INIT = 4'h8;
LUT5 lut_inst_40 (
  .F(lut_f_40),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_40.INIT = 32'h00100000;
LUT2 lut_inst_41 (
  .F(lut_f_41),
  .I0(ce),
  .I1(lut_f_40)
);
defparam lut_inst_41.INIT = 4'h8;
LUT5 lut_inst_42 (
  .F(lut_f_42),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_42.INIT = 32'h00200000;
LUT2 lut_inst_43 (
  .F(lut_f_43),
  .I0(ce),
  .I1(lut_f_42)
);
defparam lut_inst_43.INIT = 4'h8;
LUT5 lut_inst_44 (
  .F(lut_f_44),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_44.INIT = 32'h00400000;
LUT2 lut_inst_45 (
  .F(lut_f_45),
  .I0(ce),
  .I1(lut_f_44)
);
defparam lut_inst_45.INIT = 4'h8;
LUT5 lut_inst_46 (
  .F(lut_f_46),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17]),
  .I4(ad[18])
);
defparam lut_inst_46.INIT = 32'h00800000;
LUT2 lut_inst_47 (
  .F(lut_f_47),
  .I0(ce),
  .I1(lut_f_46)
);
defparam lut_inst_47.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b1;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000003FFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFC00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFE00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFE000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_19 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFF;
defparam prom_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000007FFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000003FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFC0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_32 = 256'h000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000007FFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000003FFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b1;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFF00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFFF80000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0B = 256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000003FFFFFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFFFFFFFFE000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hFFFFF000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_24 = 256'h000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam prom_inst_1.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_27 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000;
defparam prom_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000001FFFFFFF;
defparam prom_inst_1.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000FFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFC000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFC000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3A = 256'hFFFFFC000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b1;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000;
defparam prom_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFF;
defparam prom_inst_2.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_13 = 256'hFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_16 = 256'h00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_2.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_19 = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000;
defparam prom_inst_2.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFF;
defparam prom_inst_2.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000FFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFE0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2C = 256'hFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2F = 256'h000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_2.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_32 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000;
defparam prom_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000001FFFF;
defparam prom_inst_2.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFC000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b1;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_05 = 256'hFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_08 = 256'h0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_3.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0B = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
defparam prom_inst_3.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000003FFF;
defparam prom_inst_3.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFF8000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1E = 256'hFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_21 = 256'hC000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_24 = 256'h00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000;
defparam prom_inst_3.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFF;
defparam prom_inst_3.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_37 = 256'hFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3A = 256'hF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3D = 256'h000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_9),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b1;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FF;
defparam prom_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000FFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_10 = 256'hFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_13 = 256'hFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_16 = 256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
defparam prom_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000003F;
defparam prom_inst_4.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2C = 256'hFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2F = 256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000;
defparam prom_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007;
defparam prom_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFF;
defparam prom_inst_4.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_11),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b1;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_02 = 256'hFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_05 = 256'hFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_08 = 256'h00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000;
defparam prom_inst_5.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001;
defparam prom_inst_5.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFF;
defparam prom_inst_5.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000007FFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1B = 256'hFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1E = 256'hFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_21 = 256'h000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_5.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_24 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000;
defparam prom_inst_5.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFFFF;
defparam prom_inst_5.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_34 = 256'hFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_37 = 256'hFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3A = 256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam prom_inst_5.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3D = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000;
defparam prom_inst_5.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_13),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b1;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFF;
defparam prom_inst_6.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0D = 256'hFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_10 = 256'hFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_13 = 256'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam prom_inst_6.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_16 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000;
defparam prom_inst_6.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000FFFFFF;
defparam prom_inst_6.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_26 = 256'hFFFFFFFFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_29 = 256'hFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_2C = 256'h00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_6.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_2F = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000;
defparam prom_inst_6.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFF;
defparam prom_inst_6.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_15),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b1;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_02 = 256'hFFFFFFF8000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_05 = 256'h000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_7.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_08 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000;
defparam prom_inst_7.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000003FFFF;
defparam prom_inst_7.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000001FFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_11 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_12 = 256'hFFFFF00000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_15 = 256'h00000000000000000000000000000000000000000000000000000000000001FF;
defparam prom_inst_7.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_7.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000007FFFFFFFFF;
defparam prom_inst_7.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000;
defparam prom_inst_7.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1B = 256'h000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000;
defparam prom_inst_7.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1E = 256'h00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_21 = 256'h000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_24 = 256'h00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_27 = 256'h0000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_28 = 256'hFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_2A = 256'h000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_2B = 256'hFFFFF80000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_2D = 256'h0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_7.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_31 = 256'h000000000000000000000000000000000000000000000000000000000000FFFF;
defparam prom_inst_7.INIT_RAM_32 = 256'h1FFE1FFFFF9FFFFFFFF7FFFE7FBFFFFFFFF7FFE7FFFFFFFFFFFFFC0000000000;
defparam prom_inst_7.INIT_RAM_33 = 256'hFFFF7FFFFFFFFFE7FEFFFFFE7FFFFFF9FFFEFFFFE1FFFFFF7FFEFFFFFC7FFFFF;
defparam prom_inst_7.INIT_RAM_34 = 256'h00000000000000000000000000000000000000000000000000003FFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_35 = 256'h3F0003FF0003F8001F1FFFCF8FF3FFC7FCFFF9FFFFFFFE000000000000000000;
defparam prom_inst_7.INIT_RAM_36 = 256'hFF1F8003FC7FFFFC3FFFE000FFF87FFF8007FFFE3FFE7FFE0001F8001F00007E;
defparam prom_inst_7.INIT_RAM_37 = 256'hC000000000000FFFFFFFFE00000000000000000000001FFFFFFFFFFF1FFE3F3F;
defparam prom_inst_7.INIT_RAM_38 = 256'h0003F8001F1FFF8F8FE3FF83F8FFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_39 = 256'hFC7FFFFC1FFFC000FFF83FFF0003FFFE3FFC7FFE0000F0000F00007E3F0001FF;
defparam prom_inst_7.INIT_RAM_3A = 256'h00000FFFFFFFFF00000000000000000000000FFFFFFFFFFF0FFE3F1FFF0F0003;
defparam prom_inst_7.INIT_RAM_3B = 256'h0F0FFF8F87E1FF83F87FF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000;
defparam prom_inst_7.INIT_RAM_3C = 256'h1FFFC000FFF83FFF0383FFFE3FFC7FFE0001F8000F00007E3F0003FE0003F800;
defparam prom_inst_7.INIT_RAM_3D = 256'hFFFFFFC00000000000000000000001FFFFFFFFFF0FFE1F1FFF0F0003FC7FFFFC;
defparam prom_inst_7.INIT_RAM_3E = 256'h87F1FF83FC7FF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FF;
defparam prom_inst_7.INIT_RAM_3F = 256'h7FF81FFF07C0FFFE1FFC3FFFFC0FFFFE0FFC07FE1F03FFFE07E3FFFE0F87FF8F;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_17),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b1;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'h0000000000000000000000FFFFFFFFFF0FFE1F0FFF0FFFC1FC7FFFFC1FFF81F8;
defparam prom_inst_8.INIT_RAM_01 = 256'hFC7FF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFF0;
defparam prom_inst_8.INIT_RAM_02 = 256'h1FF0FFFE1FFE3FFFFC3FFFFF8FFF0FFE1F87FFFC3FE1FFFF0FC7FF8FC7F0FF81;
defparam prom_inst_8.INIT_RAM_03 = 256'h000000000000007FFFFFFFFF87FF0F8FFF0FFFE1FC7FFFFC0FFF87F87FF81FFF;
defparam prom_inst_8.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFC00000000;
defparam prom_inst_8.INIT_RAM_05 = 256'h0FFE1FFFFE3FFFFF8FFF1FFF1F87FFFC3FF1FFFF8FC7FF8FC7F0FF81FC7FF8FF;
defparam prom_inst_8.INIT_RAM_06 = 256'h0000003FFFFFFFFFC7FF0FC7FF0FFFF0FC3FFFFC07FF0FFC3FF80FFF1FF8FFFF;
defparam prom_inst_8.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFC0000000000000000;
defparam prom_inst_8.INIT_RAM_08 = 256'hFE3FFFFF8FFF0FFF1FC3FFFC3FF1FFFF8FC3FF8FC7F8FF81FC3FF8FFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_09 = 256'hFFFFFFFFC7FF8FC7FF0FFFF0FC3FFFFC07FF0FFC3FF80FFF1FF87FFF0FFE1FFF;
defparam prom_inst_8.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFF00000000000000000000000F;
defparam prom_inst_8.INIT_RAM_0B = 256'h87FF0FFF0FE1FFFC3FF0FFFF87E3FF8FC3F8FF80FC3FF87FFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0C = 256'hC7FF8FC7FF0FFFF0FE1FFFFC47FF8FFE3FF807FFBFF87FFF8FFF1FFFFE1FFFFF;
defparam prom_inst_8.INIT_RAM_0D = 256'hFFFFFFFFFC000000000003FFFFFFFFFFC00000000000000000000007FFFFFFFF;
defparam prom_inst_8.INIT_RAM_0E = 256'h0FE1FFFC3FF0FFFF87E1FF8FE3F8FF80FC3FF87FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0F = 256'hFF0FFFF8FE1FFFFC63FF8FFE3FF867FFBFFC3FFF8FFF1FFFFE1FFFFF87FF87FF;
defparam prom_inst_8.INIT_RAM_10 = 256'hFC000000000001FFFFFFFFFFC00000000000000000000003FFFFFFFFC7FF8FC3;
defparam prom_inst_8.INIT_RAM_11 = 256'h3FF0FFFFC7F1FF8FE3F8FF08FE3FFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_12 = 256'hFF1FFFFC63FF87FE3FF863FFFFFC3FFF8FFF1FFFFF1FFFFF87FF87FF0FF0FFFE;
defparam prom_inst_8.INIT_RAM_13 = 256'h000001FFFFFFFFFFE00000000000000000000001FFFFFFFFC7FF8FE1FF0FFFF8;
defparam prom_inst_8.INIT_RAM_14 = 256'hC7F1FF8FE3F8FF18FE1FFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000;
defparam prom_inst_8.INIT_RAM_15 = 256'h71FFC7FE3FF863FFFFFC3FFF8FFF1FFFFF1FFFFFC3FF87FF8FF87FFE1FF8FFFF;
defparam prom_inst_8.INIT_RAM_16 = 256'hFFFFFFFFF00000000000000000000000FFFFFFFFC3FF8FF1FF0FFFF8FF1FFFFC;
defparam prom_inst_8.INIT_RAM_17 = 256'hE1FC7F18FF1FFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000001FF;
defparam prom_inst_8.INIT_RAM_18 = 256'h3FF863FFFFFC3FFF8FFF1FFFFF1FFFFFC3FFC7FF87F87FFE1FF87FFFC3F8FF8F;
defparam prom_inst_8.INIT_RAM_19 = 256'hF800000000000000000000007FFFFFFFC3FF87F1FF0FFFF87F1FFFFC79FFC7FE;
defparam prom_inst_8.INIT_RAM_1A = 256'hFF1FFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000001FFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1B = 256'hFFFC3FFF87FF8FFFFF0FFFFFE3FFC7FF87FC3FFF1FF87FFFC3F8FF8FE1FC7F18;
defparam prom_inst_8.INIT_RAM_1C = 256'h00000000000000003FFFFFFFE3FFC7F1FF0FFFF87F1FFFFC78FFC7FE1FF871FF;
defparam prom_inst_8.INIT_RAM_1D = 256'hFFFFFFFF00000000000001F00001FFFFFE000000000000FFFFFFFFFFF8000000;
defparam prom_inst_8.INIT_RAM_1E = 256'h87FF8FFFFF8FFFFFC3FFC7FFC7FE1FFF8FF87FFFC3F87F8FF1FC7F187F1FFE3F;
defparam prom_inst_8.INIT_RAM_1F = 256'h000000001FFFFFFFE1FFC3F8FF0FFFF87F1FFFFC78FFC3FE1FF871FFFFF83FFF;
defparam prom_inst_8.INIT_RAM_20 = 256'h000000000000000000003FFFFF000000000000FFFFFFFFFFFC00000000000000;
defparam prom_inst_8.INIT_RAM_21 = 256'hFF8FFFFFC3FFC7FFC7FE1FFF83F87FFF83FC7F8FF1FC3F1C7F1FFE3FFFFFFFFC;
defparam prom_inst_8.INIT_RAM_22 = 256'h0FFFFFFFF1FFC3F87F0FFFF83F0FFFFC7C7FE0FE0FF878FFFFF07FFFC3FF8FFF;
defparam prom_inst_8.INIT_RAM_23 = 256'h0000000000001FFFFF0000000000007FFFFFFFFFFE0000000000000000000000;
defparam prom_inst_8.INIT_RAM_24 = 256'hC3FFC3FFC7FF0FFFC3F87FFF81FE3F8FF1FE3F1C7F1FFE3FFFFFFFF800000000;
defparam prom_inst_8.INIT_RAM_25 = 256'hF1FFE3FC7F0FFFF83F8FFFFC7C7FF07E0FF878FFFFE0FFFFC3FF87FFFF8FFFFF;
defparam prom_inst_8.INIT_RAM_26 = 256'h00000FFFFF0000000000007FFFFFFFFFFF000000000000000000000007FFFFFF;
defparam prom_inst_8.INIT_RAM_27 = 256'hC7FF0FFFE0F87FC001FE3F8FF0FE3E1E3F0FFE1FFFFFFFF80000000000000000;
defparam prom_inst_8.INIT_RAM_28 = 256'h7F0FFC183F87FFFC7E3FF83E0FF87C7FFFC0FFFFE3FF87FFFF87FFF041FFE3FF;
defparam prom_inst_8.INIT_RAM_29 = 256'hFF8000000000007FFFFFFFFFFF000000000000000000000003FFFFFFF1FFE3FC;
defparam prom_inst_8.INIT_RAM_2A = 256'hE0003FC001FE1F8FF8FE3E3E3F0FFE1FFFFFFFFC0000000000000000000007FF;
defparam prom_inst_8.INIT_RAM_2B = 256'h3F87FFFC7E3FF8000FF87C7FFE01FFFFE3FFC7FFFF87FFF0C1FFE3FFC3FF87FF;
defparam prom_inst_8.INIT_RAM_2C = 256'h0000003FFFFFFFFFFF800000000000000000000001FFFFFFF1FFE3FE3F0FFC18;
defparam prom_inst_8.INIT_RAM_2D = 256'h01FF1F8FF8FF1E3E3F87FF1FFFFFFFFE0000000000000000000003FFFF800000;
defparam prom_inst_8.INIT_RAM_2E = 256'h7E3FFC000FF8FE3FFC07FFFFE3FFC7FFFFC7FFF0C1FFE1FFC3FFC3FFF0003FC0;
defparam prom_inst_8.INIT_RAM_2F = 256'hFFFFFFFFFF800000000000000000000001FFFFFFF1FFE3FE1F0FFC083FC7FFFC;
defparam prom_inst_8.INIT_RAM_30 = 256'hF8FF1E3E3F87FF0FFFFFFFFE0000000000000000000003FFFF8000000000003F;
defparam prom_inst_8.INIT_RAM_31 = 256'h0FF87E3FF80FFFFFE3FFC7FFFFC3FFFFE0FFE1FFE3FFE3FFF0003FFFE1FF0F8F;
defparam prom_inst_8.INIT_RAM_32 = 256'hFFC00000000000000000000000FFFFFFF1FFE1FE1F0FFFFE3FC7FFFC7F1FFC00;
defparam prom_inst_8.INIT_RAM_33 = 256'h3FC7FF0FFFFFFFFF0000000000000000000001FFFFC000000000001FFFFFFFFF;
defparam prom_inst_8.INIT_RAM_34 = 256'hF81FFFFFE3FFE3FFFFC3FFFFE0FFF1FFE1FFE1FFE0781FFFF0FF8F8FF87F1E3E;
defparam prom_inst_8.INIT_RAM_35 = 256'h0000000000000000007FFFFFF0FFF1FF1F0FFFFE1FC7FFFC7E0FFC0F8FF87E1F;
defparam prom_inst_8.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFF0000000000001FFFFC000000000001FFFFFFFFFFFE00000;
defparam prom_inst_8.INIT_RAM_37 = 256'hE1FFE3FFFFE3FFFFF0FFF1FFF1FFF0FFE1FE1FFFF0FF8F8FF87F1C7E3FC7FF8F;
defparam prom_inst_8.INIT_RAM_38 = 256'h00000000003FFFFFF8FFF1FF8F0FFFFE1FC7FFFC1C0FF87F87F8301FF07FFFFF;
defparam prom_inst_8.INIT_RAM_39 = 256'hFFFFFFFFFC000000000000FFFFC000000000001FFFFFFFFFFFE0000000000000;
defparam prom_inst_8.INIT_RAM_3A = 256'hFFE3FFFFF8FFF1FFF1FFF8FFE3FF1FFFF0FFC78FF87F1C7E1FC7FF8FFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3B = 256'h003FFFFFF87FF0FF8F0FFFFE1FC7FFFC000FF87FC7F8000FF0FFFFFFF1FFE3FF;
defparam prom_inst_8.INIT_RAM_3C = 256'hFE000000000000FFFFE000000000000FFFFFFFFFFFE000000000000000000000;
defparam prom_inst_8.INIT_RAM_3D = 256'hF8FFF0FFF1FFF87FE3FF1FFFF8FFC38FFC7F0C7F1FC7FF8FFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3E = 256'hF87FF0FF870FFFFF0FC3FFFC0007F87FC3F8000FF0FFFFFFF0FFE3FFFFE3FFFF;
defparam prom_inst_8.INIT_RAM_3F = 256'h0000007FFFE000000000000FFFFFFFFFFFF000000000000000000000001FFFFF;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_19),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b1;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'hF1FFFC3FE3FF1FFFF87FE38FFC3F0C7F0FC7FF8FFFFFFFFFFFFFFFFFFF000000;
defparam prom_inst_9.INIT_RAM_01 = 256'hC70FFFFF0FE3FFFC1F83F87FC3F83E0FF1FFFFFFF0FFE1FFFFE3FFFFF8FFF0FF;
defparam prom_inst_9.INIT_RAM_02 = 256'hFFE000000000000FFFFFFFFFFFF000000000000000000000000FFFFFFC7FF0FF;
defparam prom_inst_9.INIT_RAM_03 = 256'hE3FF1FFFF87FE38FFE3F8C7F0FC3FF87FFFFFFFFFFFFFFFFFFC000000000007F;
defparam prom_inst_9.INIT_RAM_04 = 256'h0FE3FFFC3FC3F87FC3F83F87F1FFFFFFF8FFE1FFFFE3FFFFF87FF8FFF1FFFC3F;
defparam prom_inst_9.INIT_RAM_05 = 256'h00000007FFFFFFFFFFF800000000000000000000000FFFFFFC7FF8FFE30FFFFF;
defparam prom_inst_9.INIT_RAM_06 = 256'hFC7FE38FFE3F847F8FC3FFC7FFFFFFFFFFFFFFFFFFC000000000007FFFF00000;
defparam prom_inst_9.INIT_RAM_07 = 256'h3FE3FC7FE3F87FC7F1FFFFFFF8FFF1FFFFE1FFFFF87FF8FFF0FFFE1FE3FF0FFF;
defparam prom_inst_9.INIT_RAM_08 = 256'hFFFFFFFFFFF8000000000000000000000007FFFFFC7FF8FFE30FFFFF0FE1FFFC;
defparam prom_inst_9.INIT_RAM_09 = 256'hFE3FC47F8FE1FFC7FFFFFFFFFFFFFFFFFFE000000000003FFFF0000000000007;
defparam prom_inst_9.INIT_RAM_0A = 256'hE3F87FC3F1FFF3FFF8FFF1FFFFE1FFFFF87FF87FF0FFFF0FE1FF0FFFFC7FF00F;
defparam prom_inst_9.INIT_RAM_0B = 256'hFFF8000000000000000000000003FFFFFC7FF87FE20FFFFF8FE1FCFC7FE3FC7F;
defparam prom_inst_9.INIT_RAM_0C = 256'h8FE1FFC7FFFFFFFFFFFFFFFFFFF000000000003FFFF8000000000003FFFFFFFF;
defparam prom_inst_9.INIT_RAM_0D = 256'hF1FFF1FFF87FF0FFFFF0FFFFFC3FF87FF8FFFF0FE1FF8FFFFC7FF00FFE3FC07F;
defparam prom_inst_9.INIT_RAM_0E = 256'h00000000000000000003FFFFFC3FF87FF00FFFFF87F1FC7C7FF1FC7FE3F87FE3;
defparam prom_inst_9.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFF800000000003FFFF8000000000003FFFFFFFFFFF80000;
defparam prom_inst_9.INIT_RAM_10 = 256'hF87FF0FFFFF0FFFFFC3FF87FF87FFF87F1FF87FFFC7FF80FFE3FC07F8FF1FFC3;
defparam prom_inst_9.INIT_RAM_11 = 256'h000000000001FFFFFE3FFC7FF00FFFFF87F1FC3C7FF0FC7FE1F87FF1F0FFE1FF;
defparam prom_inst_9.INIT_RAM_12 = 256'hFFFFFFFFFFF800000000001FFFF8000000000003FFFFFFFFFFF8000000000000;
defparam prom_inst_9.INIT_RAM_13 = 256'hFFF0FFFFFC3FFC7FFC7FFFC7F1FFC7FFFC3FF80FFE1FC07F8FF1FFC3FFFFFFFF;
defparam prom_inst_9.INIT_RAM_14 = 256'h0000FFFFFE1FF87FF80FFFFF87F0FC3C7FF8FC7FF1F87FF1F8FFE1FFFC7FF0FF;
defparam prom_inst_9.INIT_RAM_15 = 256'hFFF800000000001FFFFC000000000003FFFFFFFFFFFC00000000000000000000;
defparam prom_inst_9.INIT_RAM_16 = 256'hFE3FFC3FFC7FFFC3F0FFC7FFFC3FFC0FFE1FC0FF87F07F83FFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_17 = 256'hFF0FF87FF80FFFFFC7F8FC3C7FF8FC7FF1F87FF0F87FC1FFFC1FF0FFFFF8FFFF;
defparam prom_inst_9.INIT_RAM_18 = 256'h0000000FFFFC000000000001FFFFFFFFFFFC000000000000000000000000FFFF;
defparam prom_inst_9.INIT_RAM_19 = 256'hFC7FFFC1F0FFC7FFFC1FFC0FFF0FC0FFC7F87F83FFFFFFFFFFFFFFFFFFFE0000;
defparam prom_inst_9.INIT_RAM_1A = 256'hFC0FFFFFC3F87C3C7FFC7C3FF0F87FF8FC3FC1FFFE1FE0FFFFF8FFFFFE3FFE3F;
defparam prom_inst_9.INIT_RAM_1B = 256'hFFFE000000000001FFFFFFFFFFFC0000000000000000000000007FFFFF07F87F;
defparam prom_inst_9.INIT_RAM_1C = 256'hF8FFC7FFFC1FFE0FFF0FE0FFC7F83F87FFFFFFFFFFFFFFFFFFFE00000000000F;
defparam prom_inst_9.INIT_RAM_1D = 256'h83F87C3C7FFC7C3FF0F8FFF87C3FC3FFFF0FE0FFFFF8FFFFFE3FFE3FFC7FFFC1;
defparam prom_inst_9.INIT_RAM_1E = 256'h00000000FFFFFFFFFFFC0000000000000000000000007FFFFF87F07FFC0FFFFF;
defparam prom_inst_9.INIT_RAM_1F = 256'h381FFE0FFF8FE1FFC3FC0607FFFFFFFFFFFFFFFFFFFE00000000000FFFFE0000;
defparam prom_inst_9.INIT_RAM_20 = 256'h7FFC3E3FF0F8FFFC7E0203FFFF0101FFFFF8FFFC983FFE3FFC7F8181F8FFC7FC;
defparam prom_inst_9.INIT_RAM_21 = 256'hFFFFFFFFFFFC0000000000000000000000003FFFFF81E0FFFE1FFF0183FC387C;
defparam prom_inst_9.INIT_RAM_22 = 256'hFF8FF1FFE3FE000FFFFFFFFFFFFFFFFFFFFF000000000007FFFE000000000000;
defparam prom_inst_9.INIT_RAM_23 = 256'hF8F8FFFC7F8007FFFFC003FFFFF8FFF8003FFE3FFE7F0001F8FFC7F0001FFF0F;
defparam prom_inst_9.INIT_RAM_24 = 256'hFFFE0000000000000000000000003FFFFFE000FFFE1FFE0003FE007C7FFE3E7F;
defparam prom_inst_9.INIT_RAM_25 = 256'hF3FF801FFFFFFFFFFFFFFFFFFFFF800000000007FFFE000000000000FFFFFFFF;
defparam prom_inst_9.INIT_RAM_26 = 256'h7FC00FFFFFE007FFFFFCFFF0003FFE3FFE7E0001F9FFE7F0001FFF0FFF8FF1FF;
defparam prom_inst_9.INIT_RAM_27 = 256'h000000000000000000001FFFFFF001FFFF1FFE0003FF00FC7FFF3E7FFCF9FFFE;
defparam prom_inst_9.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFF800000000003FFFF0000000000007FFFFFFFFFFE0000;
defparam prom_inst_9.INIT_RAM_29 = 256'hFFE007FFFFFDFFF8003FFF7FFEFF0001FDFFEFF8003FFF9FFFDFFBFFF7FFC01F;
defparam prom_inst_9.INIT_RAM_2A = 256'h0000000000001FFFFFF803FFFF3FFF0007FF00FEFFFF3EFFFFFFFFFFFFC00FFF;
defparam prom_inst_9.INIT_RAM_2B = 256'hFFFFFFFFFFFF800000000003FFFF0000000000007FFFFFFFFFFE000000000000;
defparam prom_inst_9.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2D = 256'h00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFBFFF;
defparam prom_inst_9.INIT_RAM_2E = 256'hFFFFC00000000003FFFF8000000000003FFFFFFFFFFE00000000000000000000;
defparam prom_inst_9.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_31 = 256'h00000003FFFF8000000000003FFFFFFFFFFE0000000000000000000000000FFF;
defparam prom_inst_9.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_9.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_34 = 256'hFFFF8000000000003FFFFFFFFFFC00000000000000000000000007FFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001;
defparam prom_inst_9.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_37 = 256'h000000003FFFFFFFFFFC00000000000000000000000007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFFC000;
defparam prom_inst_9.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_3A = 256'h1FFFFFFFFFFC00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFC00000000000;
defparam prom_inst_9.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_3D = 256'hFFFC00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFC000000000001FFFFFFF;
defparam prom_inst_9.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_21),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b1;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFF00000000000FFFFE000000000000FFFFFFFFFFC0000;
defparam prom_inst_10.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_03 = 256'h00000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_04 = 256'hFFFFFFFFFFFFF800000000007FFFE000000000000FFFFFFFFFFC000000000000;
defparam prom_inst_10.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_06 = 256'h000001FFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_07 = 256'hFFFFFC00000000007FFFE000000000000FFFFFFFFFFC00000000000000000000;
defparam prom_inst_10.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFE3C7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0A = 256'h000000003FFFF0000000000007FFFFFFFFFC00000000000000000000000001FF;
defparam prom_inst_10.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_10.INIT_RAM_0C = 256'hFFFFFFFFF10FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0D = 256'h3FFFF0000000000007FFFFFFFFF800000000000000000000000000FFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000;
defparam prom_inst_10.INIT_RAM_0F = 256'hF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_10 = 256'h0000000003FFFFFFFFF800000000000000000000000000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000003FFFF800;
defparam prom_inst_10.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_13 = 256'h03FFFFFFFFF800000000000000000000000000FFFFFFFFFFFFFFFFFFF00FFFFF;
defparam prom_inst_10.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000003FFFF80000000000;
defparam prom_inst_10.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_16 = 256'hFFF8000000000000000000000000007FFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFF8000000000003FFFFFF;
defparam prom_inst_10.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_19 = 256'h00000000000000000000007FFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFF00000000001FFFFC000000000001FFFFFFFFF00000;
defparam prom_inst_10.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1C = 256'h000000000000003FFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1D = 256'hFFFFFFFFFFFFFF00000000000FFFFC000000000001FFFFFFFFF0000000000000;
defparam prom_inst_10.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1F = 256'h0000003FFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_20 = 256'hFFFFFF00000000000FFFFC000000000001FFFFFFFFF000000000000000000000;
defparam prom_inst_10.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_23 = 256'h000000000FFFFE000000000000FFFFFFFFE0000000000000000000000000003F;
defparam prom_inst_10.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_10.INIT_RAM_25 = 256'hFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_26 = 256'h07FFFE000000000000FFFFFFFFE0000000000000000000000000003FFFFFFFFF;
defparam prom_inst_10.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000;
defparam prom_inst_10.INIT_RAM_28 = 256'hFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_29 = 256'h00000000007FFFFFFFE0000000000000000000000000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_2A = 256'hFFFFC000FFFFFFF1FFFE0003FFFFFFFFFFFFFFFFFFFFFF800000000007FFFF00;
defparam prom_inst_10.INIT_RAM_2B = 256'hF1FFE3FFFF3FFC7FFFC0003FFF80001FFFFC00FFFFFFC001FFFF0000FFFF3FFD;
defparam prom_inst_10.INIT_RAM_2C = 256'h007FFFFFFFC0000000000000000000000000001FFFC7FFFE3FF9FFFFF003FFFF;
defparam prom_inst_10.INIT_RAM_2D = 256'h7FFFFFE1FFFE0000FFFFFFFFFFFFFFFFFFFFFFC00000000007FFFF0000000000;
defparam prom_inst_10.INIT_RAM_2E = 256'hFE1FFC3FFF80001FFF00000FFFF8003FFFFF0000FFFC00007FFC0FF07FFF8000;
defparam prom_inst_10.INIT_RAM_2F = 256'hFF80000000000000000000000000000FFF83FFFC1FF0FFFFC000FFFFE0FF81FF;
defparam prom_inst_10.INIT_RAM_30 = 256'hFFFC0000FFFFFFFFFFFFFFFFFFFFFFC00000000003FFFF0000000000007FFFFF;
defparam prom_inst_10.INIT_RAM_31 = 256'hFF80001FFF00000FFFF0001FFFFE00007FFC00007FFC07F03FFF00003FFFFFE0;
defparam prom_inst_10.INIT_RAM_32 = 256'h00000000000000000000000FFF83FFF80FE07FFFC0007FFFE0FF81FFFC0FF83F;
defparam prom_inst_10.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFC00000000003FFFF0000000000007FFFFFFF800000;
defparam prom_inst_10.INIT_RAM_34 = 256'hFF00000FFFE0000FFFFE00007FFC00007FFC07F03FFF00003FFFFFE0FFFC0000;
defparam prom_inst_10.INIT_RAM_35 = 256'h000000000000000FFF83FFF80FE07FFF80003FFFE07F01FFFC0FF81FFF80001F;
defparam prom_inst_10.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFC00000000001FFFF8000000000003FFFFFFF00000000000000;
defparam prom_inst_10.INIT_RAM_37 = 256'hFFE00007FFFC00007FFC00007FFE03F03FFF00003FFFFFE0FFFE00007FFFFFFF;
defparam prom_inst_10.INIT_RAM_38 = 256'h0000000FFF81FFFC07E07FFF80001FFFE07F01FFFC0FF81FFF80001FFF00000F;
defparam prom_inst_10.INIT_RAM_39 = 256'hFFFFFFC00000000001FFFF8000000000003FFFFFFE0000000000000000000000;
defparam prom_inst_10.INIT_RAM_3A = 256'hFFFC00007FFE00007FFF01F03FFF80003FFFFFE0FFFE00007FFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_3B = 256'hFF81FFFE03F07FFF00001FFFE07F01FFFE0FF81FFFC0001FFF80000FFFE00007;
defparam prom_inst_10.INIT_RAM_3C = 256'h0000000001FFFFC000000000001FFFFFFE00000000000000000000000000000F;
defparam prom_inst_10.INIT_RAM_3D = 256'h7FFF00007FFF80F83FFFC0001FFFFFE0FFFE00007FFFFFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_10.INIT_RAM_3E = 256'h01F07FFF00E00FFFE07F00FFFE07F81FFFE0001FFFC0001FFFC03C03FFFC0000;
defparam prom_inst_10.INIT_RAM_3F = 256'h00FFFFC000000000001FFFFFFC000000000000000000000000000007FF81FFFF;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_23),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b1;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'hFFFFC0783FFFFFF01FFFFFE0FFFFFFE07FFFFFFFFFFFFFFFFFFFFFE000000000;
defparam prom_inst_11.INIT_RAM_01 = 256'h01F00FFFF07F00FFFE07FC1FFFFFF81FFFFC03FFFFC07E01FFFC03E03FFFF807;
defparam prom_inst_11.INIT_RAM_02 = 256'h00000000001FFFFFF8000000000000000000000000000007FF81FFFF80F07FFF;
defparam prom_inst_11.INIT_RAM_03 = 256'h3FFFFFF81FFFFFE0FFFFFFE07FFFFFFFFFFFFFFFFFFFFFF00000000000FFFFC0;
defparam prom_inst_11.INIT_RAM_04 = 256'hF07E00FFFE07FC0FFFFFFC0FFFFF03FFFFC0FF01FFFC0FF03FFFF81FFFFFC078;
defparam prom_inst_11.INIT_RAM_05 = 256'h000FFFFFF0000000000000000000000000000003FFC1FFFFC0707FFF03FC0FFF;
defparam prom_inst_11.INIT_RAM_06 = 256'h1FFFFFE0FFFFFFF07FFFFFFFFFFFFFFFFFFFFFF000000000007FFFE000000000;
defparam prom_inst_11.INIT_RAM_07 = 256'hFE07FC0FFFFFFC0FFFFF03FFFF80FF81FFFC1FF03FFFFC1FFFFFE0383FFFFFF8;
defparam prom_inst_11.INIT_RAM_08 = 256'hE0000000000000000000000000000003FFC1FFFFE0707FFE03FE07FFF03E00FF;
defparam prom_inst_11.INIT_RAM_09 = 256'h7FFFFFF07FFFFFFFFFFFFFFFFFFFFFF000000000007FFFE000000000000FFFFF;
defparam prom_inst_11.INIT_RAM_0A = 256'hFFFFFC0FFFFF03FFFF80FFC0FFFC1FF83FFFFC1FFFFFF0183FFFFFF81FFFFFE0;
defparam prom_inst_11.INIT_RAM_0B = 256'h000000000000000000000003FFC0FFFFE0307FFF07FE03FFF03C00FFFF07FC0F;
defparam prom_inst_11.INIT_RAM_0C = 256'h7FFFFFFFFFFFFFFFFFFFFFF800000000007FFFF0000000000007FFFFC0000000;
defparam prom_inst_11.INIT_RAM_0D = 256'hFFFF03FFFF81FFC0FFFC0FF83FFFFC1FFFFFF8083FFFFFF81FFFFFE07FFFFFF0;
defparam prom_inst_11.INIT_RAM_0E = 256'h0000000000000003FFC0FFFFF0003FFF0FFF03FFF03C007FFF07FC0FFFFFFC0F;
defparam prom_inst_11.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFF800000000007FFFF0000000000007FFFF8000000000000000;
defparam prom_inst_11.INIT_RAM_10 = 256'hFF81FFC0FFFC0FF83FFFFC0FFFFFFC003FFFFFF81FFFFFE07FFFFFF07FFFFFFF;
defparam prom_inst_11.INIT_RAM_11 = 256'h00000003FFC0FFFFF8003FFFFFFF03FFF83C007FFF03F80FFFFFFC0FFFFF03FF;
defparam prom_inst_11.INIT_RAM_12 = 256'hFFFFFFF800000000003FFFF0000000000007FFFF000000000000000000000000;
defparam prom_inst_11.INIT_RAM_13 = 256'h7FFC07F83FFFFC0FFFFFFE003FFFFFF81FFFFFE07FFFFFE07FFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_14 = 256'hFFC0FFFFFC003FFFFFFF83FFF83C007FFF00080FFFFFFC07FFFF03FFFF81FFE0;
defparam prom_inst_11.INIT_RAM_15 = 256'h00000000003FFFF0000000000003FFFC00000000000000000000000000000003;
defparam prom_inst_11.INIT_RAM_16 = 256'h3FFFFC0FFFFFFE001FFFF0001FFFFFF07FFFC0003FFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_11.INIT_RAM_17 = 256'hFC003FFFFFFF83FFF83C007FFF00000FFFF80007FFFF83FFFF81FFE07FFE03F0;
defparam prom_inst_11.INIT_RAM_18 = 256'h001FFFF8000000000003FFE000000000000000000000000000000003FFC0FFFF;
defparam prom_inst_11.INIT_RAM_19 = 256'hFFFFFE001FFFE0001FFFFFF03FFF80003FFFFFFFFFFFFFFFFFFFFFFC00000000;
defparam prom_inst_11.INIT_RAM_1A = 256'hFFFF83FFF838107FFF00000FFFF00007FFFF83FFFF81FFE07FFF00003FFFFC0F;
defparam prom_inst_11.INIT_RAM_1B = 256'h000000000001FF8000000000000000000000000000000001FFE0FFFFFC003FFF;
defparam prom_inst_11.INIT_RAM_1C = 256'h1FFFE0001FFFFFF03FFF80003FFFFFFFFFFFFFFFFFFFFFFC00000000001FFFF8;
defparam prom_inst_11.INIT_RAM_1D = 256'hF838107FFF00000FFFF00007FFFF83FFFF81FFF07FFF00001FFFFE0FFFFFFE00;
defparam prom_inst_11.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000FFE0FFFFFC001FFFFFFF83FF;
defparam prom_inst_11.INIT_RAM_1F = 256'h1FFFFFF03FFF80003FFFFFFFFFFFFFFFFFFFFFFE00000000001FFFFC00000000;
defparam prom_inst_11.INIT_RAM_20 = 256'hFF00000FFFF00007FFFF83FFFF81FFF07FFF00001FFFFE0FFFFFFE001FFFE000;
defparam prom_inst_11.INIT_RAM_21 = 256'h00000000000000000000000000000000FFE0FFFFFC001FFFFFFF81FFF838307F;
defparam prom_inst_11.INIT_RAM_22 = 256'h3FFF80003FFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFC0000000000000000;
defparam prom_inst_11.INIT_RAM_23 = 256'hFFF80007FFFF81FFFF81FFF07FFF80001FFFFE07FFFFFC001FFFE0000FFFFFF0;
defparam prom_inst_11.INIT_RAM_24 = 256'h000000000000000000000000FFE0FFFFF8001FFFFFFF81FFF830307FFF000007;
defparam prom_inst_11.INIT_RAM_25 = 256'h3FFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFC000000000000000000000000;
defparam prom_inst_11.INIT_RAM_26 = 256'hFFFF81FFFFC1FFF07FFF80001FFFFE07FFFFFC000FFFF0000FFFFFF83FFFC000;
defparam prom_inst_11.INIT_RAM_27 = 256'h0000000000000000FFE0FFFFF8001FFFFFFF81FFF820707FFF000007FFF80007;
defparam prom_inst_11.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFF000000000007FFFE00000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_29 = 256'hFFC0FFF03FFF80001FFFFE07FFFFF8000FFFF8000FFFFFF83FFFF0001FFFFFFF;
defparam prom_inst_11.INIT_RAM_2A = 256'h00000000FFE0FFFFF8001FFFFFFF81FFF820707FFF00FE07FFFC4007FFFF81FF;
defparam prom_inst_11.INIT_RAM_2B = 256'hFFFFFFFF000000000007FFFE0000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_2C = 256'h3FFF80001FFFFE07FFFFF8080FFFFFFC0FFFFFF83FFFFFF01FFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_2D = 256'hFFE07FFFF0001FFFFFFF81FFF800707FFF81FE07FFFFFF07FFFF81FFFFC0FFF0;
defparam prom_inst_11.INIT_RAM_2E = 256'h800000000007FFFF000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_2F = 256'h1FFFFF07FFFFF8080FFFFFFC0FFFFFF83FFFFFF81FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_30 = 256'hF0381FFFFFFF81FFF800F03FFF81FE07FFFFFF07FFFFC1FFFFE0FFF03FFF80F8;
defparam prom_inst_11.INIT_RAM_31 = 256'h0007FFFF000000000000000000000000000000000000000000000000FFE07FFF;
defparam prom_inst_11.INIT_RAM_32 = 256'hFFFFF01C0FFFFFFE0FFFFFF83FFFFFFC1FFFFFFFFFFFFFFFFFFFFFFF80000000;
defparam prom_inst_11.INIT_RAM_33 = 256'hE3FF81FFFC00F03FFF81FF07FFFFFF03FFFFC1FFFFE0FFF03FFF01FC1FFFFF07;
defparam prom_inst_11.INIT_RAM_34 = 256'h000000000000000000000000000000000000000000000000FFE07FFFE03C1FFF;
defparam prom_inst_11.INIT_RAM_35 = 256'h0FFFFFFE07FFFFF83FFFFFFC1FFFFFFFFFFFFFFFFFFFFFFF800000000003FFFF;
defparam prom_inst_11.INIT_RAM_36 = 256'hFC00F03FFF81FF07FFFFFF03FFFFC0FFFFE0FFF03FFF01FC0FFFFF07FFFFF03E;
defparam prom_inst_11.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000FFE07FFFE03C1FFFC3FF81FF;
defparam prom_inst_11.INIT_RAM_38 = 256'h07FFFFF83FFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFC00000000003FFFF80000000;
defparam prom_inst_11.INIT_RAM_39 = 256'hFF81FF03FFFFFF03FFFFC0FFFFE07FF07FFF01FC0FFFFF07FFFFF03E0FFFFFFE;
defparam prom_inst_11.INIT_RAM_3A = 256'h00000000000000000000000000000000FFF07FFFE07C1FFFC1FF81FFFC00F03F;
defparam prom_inst_11.INIT_RAM_3B = 256'h1FFFFFFC1FFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFF8000000000000000;
defparam prom_inst_11.INIT_RAM_3C = 256'hFFFFFF03FFFFC0FFFFE03FE07FFF83FC0FFFFF07FFFFE03E0FFFFFFF07FFFFF8;
defparam prom_inst_11.INIT_RAM_3D = 256'h000000000000000000000000FFF07FFFC07C1FFFC0FF81FFFC00F83FFFC1FF03;
defparam prom_inst_11.INIT_RAM_3E = 256'h1FFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFF8000000000001FFFFFFFFF00;
defparam prom_inst_11.INIT_RAM_3F = 256'hFFFFC0FFFFF03FE07FFF83FC0FFFFF07FFFFC07E0FFFFFFF07FFFFF81FFFFFFC;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_25),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b1;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'h0000000000000000FFF03FFFC0FC1FFFC0FF81FFFC01F81FFFC1FF03FFFFFF03;
defparam prom_inst_12.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFE00000000000FFFFC000000000000FFFFFFFFF8000000000;
defparam prom_inst_12.INIT_RAM_02 = 256'hFFF01FC07FFF83FE0FFFFF07FFFFC07E0FFFFFFC07FFFFF01FFFFFF81FFFFFFF;
defparam prom_inst_12.INIT_RAM_03 = 256'h00000000FFF03FFF80FC0FFFC07E03FFFC01F81FFFC1FF03FFFFFF03FFFFE0FF;
defparam prom_inst_12.INIT_RAM_04 = 256'hFFFFFFFFE00000000000FFFFC000000000000FFFFFFFFFF00000000000000000;
defparam prom_inst_12.INIT_RAM_05 = 256'h7FFF81FE0FFFFF03FFFFC07E07FFF00007FFE0001FFFC0001FFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_06 = 256'hFFF03FFF80FC0FFFE00003FFFE03F81FFFC1FF83FFF80003FFFFE0FFFFF80300;
defparam prom_inst_12.INIT_RAM_07 = 256'hE00000000000FFFFE000000000000FFFFFFFFFFC000000000000000000000000;
defparam prom_inst_12.INIT_RAM_08 = 256'h07FFFF03FFFFC0FE07FFE00007FFC0001FFF80001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_09 = 256'h80FC0FFFF00003FFFE03F81FFFC1FF83FFF00001FFFFE0FFFFF800007FFF81FE;
defparam prom_inst_12.INIT_RAM_0A = 256'h00007FFFE000000000000FFFFFFFFFFE000000000000000000000000FFF83FFF;
defparam prom_inst_12.INIT_RAM_0B = 256'hFFFF80FE07FFE00007FFC0000FFF80000FFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam prom_inst_12.INIT_RAM_0C = 256'hF00003FFFE03FC1FFFC1FF83FFF00001FFFFE0FFFFFC0000FFFF81FE07FFFF03;
defparam prom_inst_12.INIT_RAM_0D = 256'hE000000000000FFFFFFFFFFF800000000000000000000000FFF83FFF81FC0FFF;
defparam prom_inst_12.INIT_RAM_0E = 256'h07FFE00007FFC0000FFF80000FFFFFFFFFFFFFFFFFFFFFFFF800000000007FFF;
defparam prom_inst_12.INIT_RAM_0F = 256'hFE03FC1FFFC1FF81FFF80001FFFFE0FFFFFE0001FFFF81FE07FFFF03FFFF81FE;
defparam prom_inst_12.INIT_RAM_10 = 256'h000007FFFFFFFFFFE00000000000000000000000FFF83FFF01FE07FFF80007FF;
defparam prom_inst_12.INIT_RAM_11 = 256'h03FFC0000FFF80000FFFFFFFFFFFFFFFFFFFFFFFF800000000007FFFE0000000;
defparam prom_inst_12.INIT_RAM_12 = 256'hFFC0FF81FFF80001FFFFE0FFFFFF0001FFFF81FE07FFFF83FFFF01FF07FFE000;
defparam prom_inst_12.INIT_RAM_13 = 256'hFFFFFFFFE00000000000000000000000FFF83FFF03FE07FFFC0007FFFE03FC1F;
defparam prom_inst_12.INIT_RAM_14 = 256'h0FFFC0000FFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFF0000000000007FF;
defparam prom_inst_12.INIT_RAM_15 = 256'hFFF80001FFFFE0FFFFFF8003FFFF81FF07FFFF83FFFF01FF07FFE00007FFC000;
defparam prom_inst_12.INIT_RAM_16 = 256'hF00000000000000000000000FFF83FFE03FE07FFFE000FFFFE07FC1FFFC0FF81;
defparam prom_inst_12.INIT_RAM_17 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFF0000000000003FFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_18 = 256'hFFFFE0FFFFFF8007FFFF83FF0FFFFFC3FFFF83FF0FFFF00007FFE0001FFFC000;
defparam prom_inst_12.INIT_RAM_19 = 256'h0000000000000000FFF83FFF07FF0FFFFE001FFFFE0FFE1FFFE1FFC3FFF80001;
defparam prom_inst_12.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFC00000000003FFFF8000000000003FFFFFFFFFFF8000000;
defparam prom_inst_12.INIT_RAM_1B = 256'hFFFFF01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1C = 256'h00000000FFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1D = 256'hFFFFFFFFFC00000000001FFFF8000000000003FFFFFFFFFFFC00000000000000;
defparam prom_inst_12.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_20 = 256'hFE00000000001FFFF8000000000003FFFFFFFFFFFE0000000000000000000000;
defparam prom_inst_12.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_23 = 256'h00000FFFFC000000000001FFFFFFFFFFFF0000000000000000000000FFFFFFFF;
defparam prom_inst_12.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000;
defparam prom_inst_12.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_26 = 256'hFC000000000000FFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFF;
defparam prom_inst_12.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_29 = 256'h000000FFFFFFFFFFFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFE000000;
defparam prom_inst_12.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2C = 256'hFFFFFFFFFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFE000000000000FF;
defparam prom_inst_12.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2F = 256'hFFC000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFE000000000000FFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_32 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFF800000000003FFFE000000000000FFFFFFFFFFFFE00000;
defparam prom_inst_12.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_35 = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_36 = 256'hFFFFFFFFFF800000000003FFFF0000000000007FFFFFFFFFFFF0000000000000;
defparam prom_inst_12.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_39 = 256'hFFC00000000003FFFF0000000000007FFFFFFFFFFFF000000000000000000000;
defparam prom_inst_12.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3C = 256'h000003FFFF8000000000007FFFFFFFFFFFF000000000000000000000FFFFFFFF;
defparam prom_inst_12.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam prom_inst_12.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3F = 256'hFF8000000000003FFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFF;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_27),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b1;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FF;
defparam prom_inst_13.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_02 = 256'h0000003FFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFF800000;
defparam prom_inst_13.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_05 = 256'hFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFC000000000003F;
defparam prom_inst_13.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_08 = 256'hFFFC00000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFC000000000003FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0B = 256'h0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFF00000000000FFFFE000000000003FFFFFFFFFFFFC0000;
defparam prom_inst_13.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0E = 256'h00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0F = 256'hFFFFFFFFFFF000000000007FFFE000000000003FFFFFFFFFFFFE000000000000;
defparam prom_inst_13.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_12 = 256'hFFF000000000007FFFE000000000003FFFFFFFFFFFFE00000000000000000003;
defparam prom_inst_13.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_15 = 256'h0000003FFFF000000000003FFFFFFFFFFFFE00000000000000000003FFFFFFFF;
defparam prom_inst_13.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000;
defparam prom_inst_13.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_18 = 256'hFFF000000000003FFFFFFFFFFFFF00000000000000000003FFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_19 = 256'h3FF9FFC3F87FE3FFFC3FFE0007FFFFFFFFFFFFFFFFFFFFFFFFF800000000003F;
defparam prom_inst_13.INIT_RAM_1A = 256'h3FFFFFE1FFFFC003FFFC1FFFFC01FFFFFFC7FE3FFFFF80003F8000FF0000FFFF;
defparam prom_inst_13.INIT_RAM_1B = 256'h0000003FFFFFFFFFFFFF00000000000000000003FFFFF1FFC7F8FFF1FE0007FE;
defparam prom_inst_13.INIT_RAM_1C = 256'hF83FC1FFF81FFC0003FFFFFFFFFFFFFFFFFFFFFFFFFC00000000003FFFF00000;
defparam prom_inst_13.INIT_RAM_1D = 256'hFFFF0000FFFC0FFFF0007FFFFF83FC1FFFFF00003F0000FE00003FFE1FF0FF83;
defparam prom_inst_13.INIT_RAM_1E = 256'hFFFFFFFFFFFF00000000000000000003FFFFF0FF83F07FE0FC0003FE1FFFFF80;
defparam prom_inst_13.INIT_RAM_1F = 256'hF01FFC0001FFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFF800000000003F;
defparam prom_inst_13.INIT_RAM_20 = 256'hFFF807FFF0007FFFFF83FC0FFFFF00001F00007E00003FFC0FE07F81F01FC1FF;
defparam prom_inst_13.INIT_RAM_21 = 256'hFFFF00000000000000000003FFFFE07F83F03FC0FC0003FC1FFFFF80FFFE0000;
defparam prom_inst_13.INIT_RAM_22 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFF800000000003FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_23 = 256'hE0003FFFFF83FC0FFFFF00001F00007E00003FFC0FF07F81F80FC1FFF00FFC00;
defparam prom_inst_13.INIT_RAM_24 = 256'h0000000000000007FFFFF07F83F03FC0FC0001FC0FFFFF807FFE00007FF807FF;
defparam prom_inst_13.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFC00000000001FFFFC00000000003FFFFFFFFFFFFF0000;
defparam prom_inst_13.INIT_RAM_26 = 256'hFF83FC0FFFFF00001F80007E00003FFE0FF07F81FC07C1FFF007FC0001FFFFFF;
defparam prom_inst_13.INIT_RAM_27 = 256'h00000007FFFFF07F81F81FC0FC0001FC0FFFFF807FFE00007FF807FFE0001FFF;
defparam prom_inst_13.INIT_RAM_28 = 256'hFFFFFFFFFFFE00000000000FFFFC00000000003FFFFFFFFFFFFF800000000000;
defparam prom_inst_13.INIT_RAM_29 = 256'hFFFF80003F80003F00003FFE0FF07FC1FE03C1FFF007FE0001FFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2A = 256'hFFFFF07F81F81FC0FC0001FE0FFFFF803FFC00007FF803FFE0101FFFFF83FE0F;
defparam prom_inst_13.INIT_RAM_2B = 256'hFFFF00000000000FFFFC00000000003FFFFFFFFFFFFF80000000000000000007;
defparam prom_inst_13.INIT_RAM_2C = 256'h3F80003F80003FFE0FF03FC1FF03C0FFF007FF0001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2D = 256'hC1FC1FC0FE0001FE0FFFFF803FFC00007FF803FFE07C0FFFFF81FE07FFFF8000;
defparam prom_inst_13.INIT_RAM_2E = 256'h00000007FFFE00000000003FFFFFFFFFFFFF8000000000000000000FFFFFF07F;
defparam prom_inst_13.INIT_RAM_2F = 256'hF807FFFE0FF03FC1FF01C0FFF003FFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_13.INIT_RAM_30 = 256'hFE1F01FE07FFFF803FFC03C07FF801FFE07C0FFFFFC1FE07FFFFFC03FFFFE03F;
defparam prom_inst_13.INIT_RAM_31 = 256'hFFFE00000000003FFFFFFFFFFFFF8000000000000000000FFFFFF03FC1FC1FC0;
defparam prom_inst_13.INIT_RAM_32 = 256'h0FF03FC1FF80E0FFF003FFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFF000000000007;
defparam prom_inst_13.INIT_RAM_33 = 256'h07FFFF801FFC0FE07FF801FFE0FE0FFFFFC1FF07FFFFFE07FFFFF83FFE0FFFFE;
defparam prom_inst_13.INIT_RAM_34 = 256'h0000003FFFFFFFFFFFFF8000000000000000000FFFFFF03FC0FC0FC0FFFFC0FE;
defparam prom_inst_13.INIT_RAM_35 = 256'hFFC0E07FF001FFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFF0000;
defparam prom_inst_13.INIT_RAM_36 = 256'h1FFC0FF07FF801FFE0FF07FFFFC1FF07FFFFFF07FFFFF83FFE0FFFFE07F83FC1;
defparam prom_inst_13.INIT_RAM_37 = 256'hFFFFFFFFFFFF8000000000000000000FFFFFF83FC0FE0FC0FFFFE0FE07FFFF80;
defparam prom_inst_13.INIT_RAM_38 = 256'hF001FFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFF00000000003F;
defparam prom_inst_13.INIT_RAM_39 = 256'h7FF801FFF1FE07FFFFC0FF07FFFFFF07FFFFF81FFE0FFFFE07F83FC1FFE0007F;
defparam prom_inst_13.INIT_RAM_3A = 256'hFFFF8000000000000000000FFFFFF83FE0FE07C0FFFFE0FF07FFFF800FFE0FF0;
defparam prom_inst_13.INIT_RAM_3B = 256'hE0FFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFF00000000003FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_3C = 256'hFFFC07FFFFE0FF07FFFFFF07FFFFF81FFE0FFFFF07F83FC0FFE0007FF041FFFF;
defparam prom_inst_13.INIT_RAM_3D = 256'h000000000000001FFFFFF83FE0FF07C0FFFFE0FF07FFFF820FFE0FF07FF800FF;
defparam prom_inst_13.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFC00000000001FFFF00000000003FFFFFFFFFFFFF8000;
defparam prom_inst_13.INIT_RAM_3F = 256'hFFE0FF07FFFFFF03FFFFF81FFE0FFFFF07F83FC0FFF8007FF041FFFFE0FFFFFF;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_29),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b1;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'h0000001FFFFFF83FE0FF07C0FFFFE0FF07FFFF820FFE0FF03FF8307FFFFC07FF;
defparam prom_inst_14.INIT_RAM_01 = 256'hFFFFFFFFFFFFC00000000001FFFF80000000003FFFFFFFFFFFFF800000000000;
defparam prom_inst_14.INIT_RAM_02 = 256'hFFFFFF83FFFFF81FFE07FFFF07F83FE0FFF8007FF060FFFFC0FFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_03 = 256'hFFFFF81FE0FF07C0FFFFE0FF07FFFF820FFE0FF03FF8307FFFF807FFFFE0FF07;
defparam prom_inst_14.INIT_RAM_04 = 256'hFFFFC00000000001FFFF80000000003FFFFFFFFFFFFF0000000000000000003F;
defparam prom_inst_14.INIT_RAM_05 = 256'hFFF0001FFF07FFFF03F81FE0FFF8007FF0607FC000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_06 = 256'hE0FF03C1FF8000FF07FFFF8307FE03F03FF8307FFFC007FFFFE0FF03FFFFFF83;
defparam prom_inst_14.INIT_RAM_07 = 256'h00000001FFFF80000000003FFFFFFFFFFFFF0000000000000000003FFFFFFC1F;
defparam prom_inst_14.INIT_RAM_08 = 256'hFF07FFFF03F81FE07FFC007FF0707FC0007FFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_14.INIT_RAM_09 = 256'hFF8000FF03FFFF8303FF00003FF8307FFF0007FFFFE0FF03FFFFFF83FFE0001F;
defparam prom_inst_14.INIT_RAM_0A = 256'hFFFFC0000000003FFFFFFFFFFFFF0000000000000000003FFFFFFC1FE0FF83C1;
defparam prom_inst_14.INIT_RAM_0B = 256'h83FC1FF07FFC007FF0707F80007FFFFFFFFFFFFFFFFFFFFFFFFFE00000000000;
defparam prom_inst_14.INIT_RAM_0C = 256'h03FFFF0383FF80001FF8383FFE0007FFFFE0FF03FFFFFF83FFE0001FFF03FFFF;
defparam prom_inst_14.INIT_RAM_0D = 256'h0000003FFFFFFFFFFFFF0000000000000000003FFFFFFC1FE0FFC1C1FF00007F;
defparam prom_inst_14.INIT_RAM_0E = 256'h7FF8007FE0F07FC0007FFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFC000;
defparam prom_inst_14.INIT_RAM_0F = 256'h83FF80001FF8383FFC000FFFFFE0FF83FFFFFF83FFE0001FFF03FFFF83FC1FF0;
defparam prom_inst_14.INIT_RAM_10 = 256'hFFFFFFFFFFFE0000000000000000007FFFFFFC1FE07FC1C1FF80007F83FFFF07;
defparam prom_inst_14.INIT_RAM_11 = 256'hE0F83FC0007FFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFC0000000003F;
defparam prom_inst_14.INIT_RAM_12 = 256'h1FF83C1FF8001FFFFFE07F81FFFFFF83FFF0000FFF83FFFF83FC1FF07FF8003F;
defparam prom_inst_14.INIT_RAM_13 = 256'hFFFE0000000000000000007FFFFFFC1FE07FC1C1FF80007F83FFFF0783FF8000;
defparam prom_inst_14.INIT_RAM_14 = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFC0000000007FFFFFFFFF;
defparam prom_inst_14.INIT_RAM_15 = 256'hF8003FFFFFE07F81FFFFFF83FFF0000FFF83FFFF83FC0FF07FF8003FE0F83FC0;
defparam prom_inst_14.INIT_RAM_16 = 256'h00000000000000FFFFFFFC1FF07FC1C1FF80007F83FFFF07C1FFC0001FF03C1F;
defparam prom_inst_14.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFF800000000007FFFC0000000007FFFFFFFFFFFFE0000;
defparam prom_inst_14.INIT_RAM_18 = 256'hFFF07FC1FFFFFF83FFFC000FFF83FFFF83FE0FF07FF0003FE0781FE0007FFFFF;
defparam prom_inst_14.INIT_RAM_19 = 256'h000000FFFFFFFC1FF07FE0C1FFC0007F81FFFF03C1FFC0001FF03C1FF0007FFF;
defparam prom_inst_14.INIT_RAM_1A = 256'hFFFFFFFFFFFFF800000000003FFF8000000000FFFFFFFFFFFFFC000000000000;
defparam prom_inst_14.INIT_RAM_1B = 256'hFFFFFF81FFFFFC0FFF83FFFF81FE0FF07FF0103FE0701FFFF07FFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1C = 256'hFFFFFC0FF03FE001FFFFE03F81FFFF0380FFC0001FF01C0FF001FFFFFFF07FC1;
defparam prom_inst_14.INIT_RAM_1D = 256'hFFFFF800000000003FFF0000000000FFFFFFFFFFFFFC000000000000000001FF;
defparam prom_inst_14.INIT_RAM_1E = 256'hFFFFFE07FF83FFFFC1FE0FF07FF0301FE0001FFFF03FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1F = 256'hF83FF001FFFFF03FC1F8FF0000FF80781FF0000FF00FFFFFFFF03FC1FFFFFFC1;
defparam prom_inst_14.INIT_RAM_20 = 256'h000000001FFF0000000000FFFFFFFFFFFFFC000000000000000001FFFFFFFE0F;
defparam prom_inst_14.INIT_RAM_21 = 256'hFF83FFFFC1FE0FF07FE0381FE0000FFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_14.INIT_RAM_22 = 256'hFFFFF83FC1F0FF0000FF80FC1FF00007F01FFFFFFFF83FC1FFFFFFC1FFFFFF07;
defparam prom_inst_14.INIT_RAM_23 = 256'h0FFE0000000000FFFFFFFFFFFFF8000000000000000003FFFFFFFE0FF83FF001;
defparam prom_inst_14.INIT_RAM_24 = 256'hC1FE0FF03FE0781FE0000FFFF83FFFFFFFFFFFFFFFFFFFFFFFFFF00000000000;
defparam prom_inst_14.INIT_RAM_25 = 256'hC1F07F00007F80FC1FF00007F03FFFFFFFF83FC1FFFFFFC0FFFFFF07FF81FFFF;
defparam prom_inst_14.INIT_RAM_26 = 256'h000001FFFFFFFFFFFFF0000000000000000003FFFFFFFE07F83FF003FFFFF83F;
defparam prom_inst_14.INIT_RAM_27 = 256'h3FE07C1FE00007FFF83FFFFFFFFFFFFFFFFF0000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_28 = 256'h007F81FC0FF00007F03FE1FFFFF83FC1FFFFFFC0FFFFFF07FF81FFFFC1FE07F0;
defparam prom_inst_14.INIT_RAM_29 = 256'hFFFFFFFFFFF0000000000000000007FFFFFFFE07F83FF803FFFFF83FC1F07F00;
defparam prom_inst_14.INIT_RAM_2A = 256'hE00007FFF83FFFFFFFFFFFFFFFFF0000000000000000000000000000000003FF;
defparam prom_inst_14.INIT_RAM_2B = 256'h0FF00003F83FE0FFFFF83FC1FFFFFFE0FFFFFF07FFC1FFFFC1FE07F03FE07C1F;
defparam prom_inst_14.INIT_RAM_2C = 256'hFFE0000000000000000007FFFFFFFF07F83FF803FFFFF83FC0F07F00003F81FC;
defparam prom_inst_14.INIT_RAM_2D = 256'hF83FFFFFFFFFFFFFFFFE0000000000000000000000000000000003FFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_2E = 256'hF83FC0FFFFF81FC1FFFFFFE0FFFFFF07FFC1FFFFC0FF03F03FC0FC1FE00003FF;
defparam prom_inst_14.INIT_RAM_2F = 256'h0000000000000FFFFFFFFF07F83FFC03FFFFF83FE0F07F00003FC1FE0FE00003;
defparam prom_inst_14.INIT_RAM_30 = 256'hFFFFFFFFFFFE0000000000000000000000000000000007FFFFFFFFFFFFC00000;
defparam prom_inst_14.INIT_RAM_31 = 256'hFFF80F81FFFFFFE0FFFC0207FFC1FFC000FF01E03FC0FC1FE00003FFF81FFFFF;
defparam prom_inst_14.INIT_RAM_32 = 256'h00001FFFFFFFFF03F03FFC03FFFFF81FE0F03F00001FC1FE0FE00001F81F80FF;
defparam prom_inst_14.INIT_RAM_33 = 256'hFFFE000000000000000000000000000000000FFFFFFFFFFFFFC0000000000000;
defparam prom_inst_14.INIT_RAM_34 = 256'hFFFFFFE0FFF80007FFC0FF0000FF80C03F80FC1FE07F03FFF81FFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_35 = 256'hFFFFFF01E03FFC03FFE0001FE0703E03F81FC0FE07E03F81FC0F00FFFFFC0701;
defparam prom_inst_14.INIT_RAM_36 = 256'h00000000000000000000000000001FFFFFFFFFFFFF8000000000000000003FFF;
defparam prom_inst_14.INIT_RAM_37 = 256'hFFF00007FFC0FF0000FF80003F80FC0FE0FF83FFFC1FFFFFFFFFFFFFFFFE0000;
defparam prom_inst_14.INIT_RAM_38 = 256'h003FFE03FFC0001FE0203E07FC1FC0FF07E07FC0FC0700FFFFFE0001FFFFFFE0;
defparam prom_inst_14.INIT_RAM_39 = 256'h000000000000000000003FFFFFFFFFFFFF0000000000000000003FFFFFFFFF80;
defparam prom_inst_14.INIT_RAM_3A = 256'hFFE0FF0000FF80007F81FC0FE0FF81FFFC1FFFFFFFFFFFFFFFFF000000000000;
defparam prom_inst_14.INIT_RAM_3B = 256'hFFC0001FE0003E07FC0FC0FF07E07FC0FC0001FFFFFE0001FFFFFFE0FFF00003;
defparam prom_inst_14.INIT_RAM_3C = 256'h00FFFFFFFFFFFFFFFFFFFFFFFE0000000000000000007FFFFFFFFF80003FFE03;
defparam prom_inst_14.INIT_RAM_3D = 256'h007FC0007F81FE0FE0FFC0FFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000;
defparam prom_inst_14.INIT_RAM_3E = 256'hF0007E07FC0FC0FF07E07FE0FE0001FFFFFF0001FFFFFFE07FF80003FFE0FF00;
defparam prom_inst_14.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFC000000000000000000FFFFFFFFFFC0003FFE03FFC0001F;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_31),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b1;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'h7F83FE0FE0FFC0FFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFF;
defparam prom_inst_15.INIT_RAM_01 = 256'hFE07C0FF07E07FE07F0003FFFFFF0003FFFFFFE07FF80003FFE0FF00007FE000;
defparam prom_inst_15.INIT_RAM_02 = 256'hFFFFFFFFF8000000000000000001FFFFFFFFFFE0007FFF03FFC0000FF8007E07;
defparam prom_inst_15.INIT_RAM_03 = 256'hE0FFE0FFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_04 = 256'h07E0FFE07F0003FFFFFF8003FFFFFFF0FFF80003FFE0FF80007FF000FF83FE0F;
defparam prom_inst_15.INIT_RAM_05 = 256'hE0000000000000000003FFFFFFFFFFE000FFFF03FFC0000FF8007E0FFE07E0FF;
defparam prom_inst_15.INIT_RAM_06 = 256'hFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_07 = 256'hFF8007FFFFFFC007FFFFFFF0FFF80007FFF0FF8000FFF801FF83FF1FF1FFE1FF;
defparam prom_inst_15.INIT_RAM_08 = 256'h000000000007FFFFFFFFFFF000FFFF87FFE0001FFC00FF0FFF0FE1FF87F0FFF0;
defparam prom_inst_15.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFFFFFFFFFFFFFFFFFFFF80000000;
defparam prom_inst_15.INIT_RAM_0A = 256'hFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0B = 256'h000FFFFFFFFFFFFE03FFFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFFF01FFF;
defparam prom_inst_15.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFF0000000000000000;
defparam prom_inst_15.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0E = 256'hFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0F = 256'hFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFFF80000000000000000001FFFFF;
defparam prom_inst_15.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_12 = 256'h0000000000000000000C0000000000000000000000000000007FFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_15.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_15 = 256'h000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000;
defparam prom_inst_15.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_18 = 256'h0000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000;
defparam prom_inst_15.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1B = 256'h00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1E = 256'h00000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_21 = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000000001;
defparam prom_inst_15.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_28 = 256'hFFFFFFFC00000000000000000000000000000000000000000000000FFFFFFFFF;
defparam prom_inst_15.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_15.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2E = 256'h00000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000;
defparam prom_inst_15.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_31 = 256'h00000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000;
defparam prom_inst_15.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_16 (
    .DO({prom_inst_16_dout_w[30:0],prom_inst_16_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_16.READ_MODE = 1'b1;
defparam prom_inst_16.BIT_WIDTH = 1;
defparam prom_inst_16.RESET_MODE = "SYNC";
defparam prom_inst_16.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_01 = 256'hFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_04 = 256'h800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_07 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000;
defparam prom_inst_16.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFF;
defparam prom_inst_16.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1A = 256'hFFFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1D = 256'hF000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_20 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam prom_inst_16.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFF;
defparam prom_inst_16.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_33 = 256'hFFFFFFFFFE00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_36 = 256'hFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_39 = 256'h00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
defparam prom_inst_16.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FF;
defparam prom_inst_16.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_17 (
    .DO({prom_inst_17_dout_w[30:0],prom_inst_17_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_35),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_17.READ_MODE = 1'b1;
defparam prom_inst_17.BIT_WIDTH = 1;
defparam prom_inst_17.RESET_MODE = "SYNC";
defparam prom_inst_17.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF800000000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0C = 256'hFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0F = 256'hFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_12 = 256'h000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam prom_inst_17.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FF;
defparam prom_inst_17.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_25 = 256'hFFFFFFFFFFF800000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_28 = 256'hFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2B = 256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000;
defparam prom_inst_17.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000003F;
defparam prom_inst_17.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFF;
defparam prom_inst_17.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3E = 256'hFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_18 (
    .DO({prom_inst_18_dout_w[30:0],prom_inst_18_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_37),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_18.READ_MODE = 1'b1;
defparam prom_inst_18.BIT_WIDTH = 1;
defparam prom_inst_18.RESET_MODE = "SYNC";
defparam prom_inst_18.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_01 = 256'hFFFF000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_04 = 256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_18.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000007;
defparam prom_inst_18.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFF;
defparam prom_inst_18.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_17 = 256'hFFFFFFFFFFFFE00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1A = 256'hFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1D = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_18.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000;
defparam prom_inst_18.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFFFFF;
defparam prom_inst_18.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_30 = 256'hFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_33 = 256'hFFFFFC00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_36 = 256'h000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_18.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_39 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000;
defparam prom_inst_18.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFF;
defparam prom_inst_18.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_19 (
    .DO({prom_inst_19_dout_w[30:0],prom_inst_19_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_39),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_19.READ_MODE = 1'b1;
defparam prom_inst_19.BIT_WIDTH = 1;
defparam prom_inst_19.RESET_MODE = "SYNC";
defparam prom_inst_19.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_09 = 256'hFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0C = 256'hFFFFFF000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0F = 256'h0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam prom_inst_19.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_12 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000;
defparam prom_inst_19.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000003FFFFFF;
defparam prom_inst_19.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_25 = 256'hFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_28 = 256'h00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_19.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2B = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000;
defparam prom_inst_19.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFF;
defparam prom_inst_19.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3E = 256'hFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_20 (
    .DO({prom_inst_20_dout_w[30:0],prom_inst_20_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_41),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_20.READ_MODE = 1'b1;
defparam prom_inst_20.BIT_WIDTH = 1;
defparam prom_inst_20.RESET_MODE = "SYNC";
defparam prom_inst_20.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_01 = 256'h00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_20.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_04 = 256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000;
defparam prom_inst_20.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFF;
defparam prom_inst_20.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF800000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_17 = 256'hFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1A = 256'hC00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1D = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000;
defparam prom_inst_20.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFF;
defparam prom_inst_20.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFF800000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_30 = 256'hFFFFFFFFF800000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_33 = 256'hF800000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_36 = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000;
defparam prom_inst_20.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000003FFF;
defparam prom_inst_20.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000003FFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_21 (
    .DO({prom_inst_21_dout_w[30:0],prom_inst_21_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_43),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_21.READ_MODE = 1'b1;
defparam prom_inst_21.BIT_WIDTH = 1;
defparam prom_inst_21.RESET_MODE = "SYNC";
defparam prom_inst_21.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFF00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_09 = 256'hFFFFFFFFFF80000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0C = 256'hFF80000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0F = 256'h000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000;
defparam prom_inst_21.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000007FF;
defparam prom_inst_21.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000003FFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFF00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_22 = 256'hFFFFFFFFFFF80000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_25 = 256'hFFF80000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_28 = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000;
defparam prom_inst_21.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000FF;
defparam prom_inst_21.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000FFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFF80000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3B = 256'hFFFFFFFFFFFF80000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3E = 256'hFFFFC0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_22 (
    .DO({prom_inst_22_dout_w[30:0],prom_inst_22_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_45),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_22.READ_MODE = 1'b1;
defparam prom_inst_22.BIT_WIDTH = 1;
defparam prom_inst_22.RESET_MODE = "SYNC";
defparam prom_inst_22.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_01 = 256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_22.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000001F;
defparam prom_inst_22.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFFF;
defparam prom_inst_22.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000FFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_14 = 256'hFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_17 = 256'hFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1A = 256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_22.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000003;
defparam prom_inst_22.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFF;
defparam prom_inst_22.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000001FFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFF800000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFF800000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_30 = 256'hFFFFFFFE00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_33 = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_36 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000;
defparam prom_inst_22.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000007FFFFFFF;
defparam prom_inst_22.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_23 (
    .DO({prom_inst_23_dout_w[30:0],prom_inst_23_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_47),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_23.READ_MODE = 1'b1;
defparam prom_inst_23.BIT_WIDTH = 1;
defparam prom_inst_23.RESET_MODE = "SYNC";
defparam prom_inst_23.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000003FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF80000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_09 = 256'hFFFFFFFFFF8000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0C = 256'hFFC000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0F = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000;
defparam prom_inst_23.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003FFFFFFF;
defparam prom_inst_23.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[18]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[17]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_5 (
  .Q(dff_q_5),
  .D(dff_q_4),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_6 (
  .Q(dff_q_6),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_7 (
  .Q(dff_q_7),
  .D(dff_q_6),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_8 (
  .Q(dff_q_8),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_9 (
  .Q(dff_q_9),
  .D(dff_q_8),
  .CLK(clk),
  .CE(oce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(prom_inst_4_dout[0]),
  .I1(prom_inst_5_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(prom_inst_6_dout[0]),
  .I1(prom_inst_7_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(prom_inst_8_dout[0]),
  .I1(prom_inst_9_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(prom_inst_10_dout[0]),
  .I1(prom_inst_11_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(prom_inst_12_dout[0]),
  .I1(prom_inst_13_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(prom_inst_14_dout[0]),
  .I1(prom_inst_15_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(prom_inst_16_dout[0]),
  .I1(prom_inst_17_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(prom_inst_18_dout[0]),
  .I1(prom_inst_19_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(prom_inst_20_dout[0]),
  .I1(prom_inst_21_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(prom_inst_22_dout[0]),
  .I1(prom_inst_23_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_7)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_7)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_7)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_7)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_7)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_7)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_5)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_5)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_5)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_3)
);
MUX2 mux_inst_23 (
  .O(dout[0]),
  .I0(mux_o_21),
  .I1(mux_o_20),
  .S0(dff_q_1)
);
endmodule //Gowin_pROM
