//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Sun Aug 06 17:57:16 2023

module Gowin_pROM2 (dout, clk, oce, ce, reset, ad);//colorful etf

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [15:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire [26:0] promx9_inst_0_dout_w;
wire [8:0] promx9_inst_0_dout;
wire [26:0] promx9_inst_1_dout_w;
wire [8:0] promx9_inst_1_dout;
wire [26:0] promx9_inst_2_dout_w;
wire [8:0] promx9_inst_2_dout;
wire [26:0] promx9_inst_3_dout_w;
wire [8:0] promx9_inst_3_dout;
wire [26:0] promx9_inst_4_dout_w;
wire [8:0] promx9_inst_4_dout;
wire [26:0] promx9_inst_5_dout_w;
wire [8:0] promx9_inst_5_dout;
wire [26:0] promx9_inst_6_dout_w;
wire [8:0] promx9_inst_6_dout;
wire [26:0] promx9_inst_7_dout_w;
wire [8:0] promx9_inst_7_dout;
wire [26:0] promx9_inst_8_dout_w;
wire [8:0] promx9_inst_8_dout;
wire [26:0] promx9_inst_9_dout_w;
wire [8:0] promx9_inst_9_dout;
wire [26:0] promx9_inst_10_dout_w;
wire [8:0] promx9_inst_10_dout;
wire [26:0] promx9_inst_11_dout_w;
wire [8:0] promx9_inst_11_dout;
wire [26:0] promx9_inst_12_dout_w;
wire [8:0] promx9_inst_12_dout;
wire [26:0] promx9_inst_13_dout_w;
wire [8:0] promx9_inst_13_dout;
wire [26:0] promx9_inst_14_dout_w;
wire [8:0] promx9_inst_14_dout;
wire [26:0] promx9_inst_15_dout_w;
wire [8:0] promx9_inst_15_dout;
wire [30:0] prom_inst_16_dout_w;
wire [9:9] prom_inst_16_dout;
wire [30:0] prom_inst_17_dout_w;
wire [9:9] prom_inst_17_dout;
wire [30:0] prom_inst_18_dout_w;
wire [10:10] prom_inst_18_dout;
wire [30:0] prom_inst_19_dout_w;
wire [10:10] prom_inst_19_dout;
wire [30:0] prom_inst_20_dout_w;
wire [11:11] prom_inst_20_dout;
wire [30:0] prom_inst_21_dout_w;
wire [11:11] prom_inst_21_dout;
wire [30:0] prom_inst_22_dout_w;
wire [12:12] prom_inst_22_dout;
wire [30:0] prom_inst_23_dout_w;
wire [12:12] prom_inst_23_dout;
wire [30:0] prom_inst_24_dout_w;
wire [13:13] prom_inst_24_dout;
wire [30:0] prom_inst_25_dout_w;
wire [13:13] prom_inst_25_dout;
wire [30:0] prom_inst_26_dout_w;
wire [14:14] prom_inst_26_dout;
wire [30:0] prom_inst_27_dout_w;
wire [14:14] prom_inst_27_dout;
wire [30:0] prom_inst_28_dout_w;
wire [15:15] prom_inst_28_dout;
wire [30:0] prom_inst_29_dout_w;
wire [15:15] prom_inst_29_dout;
wire [26:0] promx9_inst_30_dout_w;
wire [8:0] promx9_inst_30_dout;
wire [26:0] promx9_inst_31_dout_w;
wire [8:0] promx9_inst_31_dout;
wire [26:0] promx9_inst_32_dout_w;
wire [8:0] promx9_inst_32_dout;
wire [26:0] promx9_inst_33_dout_w;
wire [8:0] promx9_inst_33_dout;
wire [26:0] promx9_inst_34_dout_w;
wire [8:0] promx9_inst_34_dout;
wire [26:0] promx9_inst_35_dout_w;
wire [8:0] promx9_inst_35_dout;
wire [26:0] promx9_inst_36_dout_w;
wire [8:0] promx9_inst_36_dout;
wire [26:0] promx9_inst_37_dout_w;
wire [8:0] promx9_inst_37_dout;
wire [30:0] prom_inst_38_dout_w;
wire [9:9] prom_inst_38_dout;
wire [30:0] prom_inst_39_dout_w;
wire [10:10] prom_inst_39_dout;
wire [30:0] prom_inst_40_dout_w;
wire [11:11] prom_inst_40_dout;
wire [30:0] prom_inst_41_dout_w;
wire [12:12] prom_inst_41_dout;
wire [30:0] prom_inst_42_dout_w;
wire [13:13] prom_inst_42_dout;
wire [30:0] prom_inst_43_dout_w;
wire [14:14] prom_inst_43_dout;
wire [30:0] prom_inst_44_dout_w;
wire [15:15] prom_inst_44_dout;
wire [15:0] prom_inst_45_dout_w;
wire [15:0] prom_inst_45_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire dff_q_7;
wire dff_q_8;
wire dff_q_9;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_49;
wire mux_o_50;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_101;
wire mux_o_102;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_153;
wire mux_o_154;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_205;
wire mux_o_206;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_257;
wire mux_o_258;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_309;
wire mux_o_310;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_361;
wire mux_o_362;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_413;
wire mux_o_414;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire mux_o_447;
wire mux_o_448;
wire mux_o_449;
wire mux_o_450;
wire mux_o_451;
wire mux_o_452;
wire mux_o_454;
wire mux_o_455;
wire mux_o_456;
wire mux_o_457;
wire mux_o_458;
wire mux_o_459;
wire mux_o_461;
wire mux_o_462;
wire mux_o_463;
wire mux_o_465;
wire mux_o_466;
wire mux_o_484;
wire mux_o_485;
wire mux_o_503;
wire mux_o_504;
wire mux_o_522;
wire mux_o_523;
wire mux_o_541;
wire mux_o_542;
wire mux_o_560;
wire mux_o_561;
wire mux_o_579;
wire mux_o_580;
wire mux_o_598;
wire mux_o_599;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT5 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_0.INIT = 32'h00000001;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(lut_f_0)
);
defparam lut_inst_1.INIT = 4'h8;
LUT5 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_2.INIT = 32'h00000002;
LUT2 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(lut_f_2)
);
defparam lut_inst_3.INIT = 4'h8;
LUT5 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_4.INIT = 32'h00000004;
LUT2 lut_inst_5 (
  .F(lut_f_5),
  .I0(ce),
  .I1(lut_f_4)
);
defparam lut_inst_5.INIT = 4'h8;
LUT5 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_6.INIT = 32'h00000008;
LUT2 lut_inst_7 (
  .F(lut_f_7),
  .I0(ce),
  .I1(lut_f_6)
);
defparam lut_inst_7.INIT = 4'h8;
LUT5 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_8.INIT = 32'h00000010;
LUT2 lut_inst_9 (
  .F(lut_f_9),
  .I0(ce),
  .I1(lut_f_8)
);
defparam lut_inst_9.INIT = 4'h8;
LUT5 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_10.INIT = 32'h00000020;
LUT2 lut_inst_11 (
  .F(lut_f_11),
  .I0(ce),
  .I1(lut_f_10)
);
defparam lut_inst_11.INIT = 4'h8;
LUT5 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_12.INIT = 32'h00000040;
LUT2 lut_inst_13 (
  .F(lut_f_13),
  .I0(ce),
  .I1(lut_f_12)
);
defparam lut_inst_13.INIT = 4'h8;
LUT5 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_14.INIT = 32'h00000080;
LUT2 lut_inst_15 (
  .F(lut_f_15),
  .I0(ce),
  .I1(lut_f_14)
);
defparam lut_inst_15.INIT = 4'h8;
LUT5 lut_inst_16 (
  .F(lut_f_16),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_16.INIT = 32'h00000100;
LUT2 lut_inst_17 (
  .F(lut_f_17),
  .I0(ce),
  .I1(lut_f_16)
);
defparam lut_inst_17.INIT = 4'h8;
LUT5 lut_inst_18 (
  .F(lut_f_18),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_18.INIT = 32'h00000200;
LUT2 lut_inst_19 (
  .F(lut_f_19),
  .I0(ce),
  .I1(lut_f_18)
);
defparam lut_inst_19.INIT = 4'h8;
LUT5 lut_inst_20 (
  .F(lut_f_20),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_20.INIT = 32'h00000400;
LUT2 lut_inst_21 (
  .F(lut_f_21),
  .I0(ce),
  .I1(lut_f_20)
);
defparam lut_inst_21.INIT = 4'h8;
LUT5 lut_inst_22 (
  .F(lut_f_22),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_22.INIT = 32'h00000800;
LUT2 lut_inst_23 (
  .F(lut_f_23),
  .I0(ce),
  .I1(lut_f_22)
);
defparam lut_inst_23.INIT = 4'h8;
LUT5 lut_inst_24 (
  .F(lut_f_24),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_24.INIT = 32'h00001000;
LUT2 lut_inst_25 (
  .F(lut_f_25),
  .I0(ce),
  .I1(lut_f_24)
);
defparam lut_inst_25.INIT = 4'h8;
LUT5 lut_inst_26 (
  .F(lut_f_26),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_26.INIT = 32'h00002000;
LUT2 lut_inst_27 (
  .F(lut_f_27),
  .I0(ce),
  .I1(lut_f_26)
);
defparam lut_inst_27.INIT = 4'h8;
LUT5 lut_inst_28 (
  .F(lut_f_28),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_28.INIT = 32'h00004000;
LUT2 lut_inst_29 (
  .F(lut_f_29),
  .I0(ce),
  .I1(lut_f_28)
);
defparam lut_inst_29.INIT = 4'h8;
LUT5 lut_inst_30 (
  .F(lut_f_30),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_30.INIT = 32'h00008000;
LUT2 lut_inst_31 (
  .F(lut_f_31),
  .I0(ce),
  .I1(lut_f_30)
);
defparam lut_inst_31.INIT = 4'h8;
LUT3 lut_inst_32 (
  .F(lut_f_32),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_32.INIT = 8'h02;
LUT3 lut_inst_33 (
  .F(lut_f_33),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_33.INIT = 8'h08;
LUT5 lut_inst_34 (
  .F(lut_f_34),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_34.INIT = 32'h00010000;
LUT2 lut_inst_35 (
  .F(lut_f_35),
  .I0(ce),
  .I1(lut_f_34)
);
defparam lut_inst_35.INIT = 4'h8;
LUT5 lut_inst_36 (
  .F(lut_f_36),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_36.INIT = 32'h00020000;
LUT2 lut_inst_37 (
  .F(lut_f_37),
  .I0(ce),
  .I1(lut_f_36)
);
defparam lut_inst_37.INIT = 4'h8;
LUT5 lut_inst_38 (
  .F(lut_f_38),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_38.INIT = 32'h00040000;
LUT2 lut_inst_39 (
  .F(lut_f_39),
  .I0(ce),
  .I1(lut_f_38)
);
defparam lut_inst_39.INIT = 4'h8;
LUT5 lut_inst_40 (
  .F(lut_f_40),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_40.INIT = 32'h00080000;
LUT2 lut_inst_41 (
  .F(lut_f_41),
  .I0(ce),
  .I1(lut_f_40)
);
defparam lut_inst_41.INIT = 4'h8;
LUT5 lut_inst_42 (
  .F(lut_f_42),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_42.INIT = 32'h00100000;
LUT2 lut_inst_43 (
  .F(lut_f_43),
  .I0(ce),
  .I1(lut_f_42)
);
defparam lut_inst_43.INIT = 4'h8;
LUT5 lut_inst_44 (
  .F(lut_f_44),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_44.INIT = 32'h00200000;
LUT2 lut_inst_45 (
  .F(lut_f_45),
  .I0(ce),
  .I1(lut_f_44)
);
defparam lut_inst_45.INIT = 4'h8;
LUT5 lut_inst_46 (
  .F(lut_f_46),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_46.INIT = 32'h00400000;
LUT2 lut_inst_47 (
  .F(lut_f_47),
  .I0(ce),
  .I1(lut_f_46)
);
defparam lut_inst_47.INIT = 4'h8;
LUT5 lut_inst_48 (
  .F(lut_f_48),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14]),
  .I4(ad[15])
);
defparam lut_inst_48.INIT = 32'h00800000;
LUT2 lut_inst_49 (
  .F(lut_f_49),
  .I0(ce),
  .I1(lut_f_48)
);
defparam lut_inst_49.INIT = 4'h8;
LUT3 lut_inst_50 (
  .F(lut_f_50),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_50.INIT = 8'h20;
LUT6 lut_inst_51 (
  .F(lut_f_51),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14]),
  .I5(ad[15])
);
defparam lut_inst_51.INIT = 64'h0001000000000000;
LUT2 lut_inst_52 (
  .F(lut_f_52),
  .I0(ce),
  .I1(lut_f_51)
);
defparam lut_inst_52.INIT = 4'h8;
pROMX9 promx9_inst_0 (
    .DO({promx9_inst_0_dout_w[26:0],promx9_inst_0_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_0.READ_MODE = 1'b1;
defparam promx9_inst_0.BIT_WIDTH = 9;
defparam promx9_inst_0.RESET_MODE = "SYNC";
defparam promx9_inst_0.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_02 = 288'h4DA6D36DCCE1F6FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF71B69B;
defparam promx9_inst_0.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_0B = 288'hFF975369B4DA6D36BB6DC6EF9FD8F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_14 = 288'hFFFFFFFFFFFBF9769B4DA6D369B4DA6CF6DBCE27B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFDFE789B4DA6D369B4DA6D36BB3DC713B7FFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA9B4DA6D369B4DA6D369B4DA6CF7FCEFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_2E = 288'hFEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDBCBB4DA6D369B4DA6D369B4DA6D36BB;
defparam promx9_inst_0.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_37 = 288'h4DA6D369B6E177FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3F1C4DA6D369B4DA6D369B;
defparam promx9_inst_0.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_0.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_1 (
    .DO({promx9_inst_1_dout_w[26:0],promx9_inst_1_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_1.READ_MODE = 1'b1;
defparam promx9_inst_1.BIT_WIDTH = 9;
defparam promx9_inst_1.RESET_MODE = "SYNC";
defparam promx9_inst_1.INIT_RAM_00 = 288'h4DA6D369B4DA6D369B4DBF1BDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDC3DA6D369B;
defparam promx9_inst_1.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_09 = 288'h3DA6D369B4DA6D369B4DA6D369B4D9EDF97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFE;
defparam promx9_inst_1.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_12 = 288'hFFFFFFFFF6DA6D369B4DA6D369B4DA6D369B4DA6D37BCEFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFF2E9ED369B4DA6D369B4DA6D369B4DA6D36DB5F7FFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFAF2ED369B4DA6D369B4DA6D369B4DAED369BBE6FFFFFF;
defparam promx9_inst_1.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_2C = 288'h4DAFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFD71369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_1.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_35 = 288'h4DA6D369B4DBF37FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF97536BB4DA6D369B4DA6D369B;
defparam promx9_inst_1.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_3E = 288'h4DA6D369B4DA6D369B4D9EC3BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_1.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC79B69B4DA6D369B;

pROMX9 promx9_inst_2 (
    .DO({promx9_inst_2_dout_w[26:0],promx9_inst_2_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_2.READ_MODE = 1'b1;
defparam promx9_inst_2.BIT_WIDTH = 9;
defparam promx9_inst_2.RESET_MODE = "SYNC";
defparam promx9_inst_2.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_07 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6E795EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFEF89B;
defparam promx9_inst_2.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_10 = 288'hFFFFC7A9B4DA6D369B4DA6D369B4DA6D369B4DA6D765DFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_19 = 288'hFFFFFFFFFFFFFE7C9B4DA6D369B4DA6D369B4DA6D369B4DA6D377CCFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFEDB4DA6D369B4DA6D369B4DA6D369B4DA6D36BB7F7FFFFFF;
defparam promx9_inst_2.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_2A = 288'hDE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7D3DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_2.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_33 = 288'h4DA6D369B6DDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9E6DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_2.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_3C = 288'h4DA6D369B4DA6D369B4D8F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDE26D369B4DA6D369B;
defparam promx9_inst_2.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_2.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_3 (
    .DO({promx9_inst_3_dout_w[26:0],promx9_inst_3_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_3.READ_MODE = 1'b1;
defparam promx9_inst_3.BIT_WIDTH = 9;
defparam promx9_inst_3.RESET_MODE = "SYNC";
defparam promx9_inst_3.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_05 = 288'h4DA6D369B4DA6D369B4DA6D369B4DAEFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6F26D369B;
defparam promx9_inst_3.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_0E = 288'hBFC71369B4DA6D369B4DA6D369B4DA6D369B4DA6DBDFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_17 = 288'hFFFFFFFFFEFF75369B4DA6D369B4DA6D369B4DA6D369B4DA6FBBFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFAF9769B4DA6D369B4DA6D369B4DA6D369B4DAEE797FFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE389B4DA6D369B4DA6D369B4DA6D369B4DA6D76DE;
defparam promx9_inst_3.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_31 = 288'h4DA6D361DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF789B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_3.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_3A = 288'h4DA6D369B4DA6D373CDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDBC7B4DA6D369B4DA6D369B;
defparam promx9_inst_3.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_3.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_4 (
    .DO({promx9_inst_4_dout_w[26:0],promx9_inst_4_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_9),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_4.READ_MODE = 1'b1;
defparam promx9_inst_4.BIT_WIDTH = 9;
defparam promx9_inst_4.RESET_MODE = "SYNC";
defparam promx9_inst_4.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_03 = 288'h4DA6D369B4DA6D369B4DA6D36BB8F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F1C4DA6D369B;
defparam promx9_inst_4.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_0C = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D367BFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1D;
defparam promx9_inst_4.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_15 = 288'hFFFFFFF5E5DA6D369B4DA6D369B4DA6D369B4DA6D369B6DEFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFDFAE26D369B4DA6D369B4DA6D369B4DA6D369B3DB7BFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFF2EA6D369B4DA6D369B4DA6D369B4DA6D369B3DEF3FFFF;
defparam promx9_inst_4.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_2F = 288'h4DBF2BDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F3ED369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_4.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_38 = 288'h4DA6D369B5DA6D3BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFDF1369B4DA6D369B4DA6D369B;
defparam promx9_inst_4.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_4.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_5 (
    .DO({promx9_inst_5_dout_w[26:0],promx9_inst_5_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_11),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_5.READ_MODE = 1'b1;
defparam promx9_inst_5.BIT_WIDTH = 9;
defparam promx9_inst_5.RESET_MODE = "SYNC";
defparam promx9_inst_5.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_01 = 288'h4DA6D369B4DA6D369B4DA6F79DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F5369B4DA6D369B;
defparam promx9_inst_5.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_0A = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6E395FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD79369B;
defparam promx9_inst_5.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_13 = 288'hFFF7EB89B4DA6D369B4DA6D369B4DA6D369B4DA6D76BEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_1C = 288'hFFFFFFFFFFFFFD3A7B4DA6D369B4DA6D369B4DA6D369B4DA6D37BCFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFF3EBB4DA6D369B4DA6D369B4DA6D369B4DA6D36DBCFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_2D = 288'h4F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDC4DA6D369B4DA6D369B4DA6D369B4DA6D367B;
defparam promx9_inst_5.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_36 = 288'h4DA6D369B9E7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFE4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_5.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_5.INIT_RAM_3F = 288'h4DA6D369B4DA6D369B4DC7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_6 (
    .DO({promx9_inst_6_dout_w[26:0],promx9_inst_6_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_13),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_6.READ_MODE = 1'b1;
defparam promx9_inst_6.BIT_WIDTH = 9;
defparam promx9_inst_6.RESET_MODE = "SYNC";
defparam promx9_inst_6.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9E9E26D369B4DA6D369B;
defparam promx9_inst_6.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_08 = 288'h4DA6D369B4DA6D369B4DA6D369B3D8F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEA6D369B;
defparam promx9_inst_6.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_11 = 288'h5F2ED369B4DA6D369B4DA6D369B4DA6D369B4DD737FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_1A = 288'hFFFFFFFFFCFBF1769B4DA6D369B4DA6D369B4DA6D369B4DB71FDFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFF75369B4DA6D369B4DA6D369B4DA6D369B4DA6C7BDFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF8F69B4DA6D369B4DA6D369B4DA6D369B4DA6EF9BF;
defparam promx9_inst_6.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_34 = 288'h4DA6DB73EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7DB89B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_6.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_3D = 288'h4DA6D369B4DAECF63DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_6.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7A7B4DA6D369B4DA6D369B;
defparam promx9_inst_6.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_7 (
    .DO({promx9_inst_7_dout_w[26:0],promx9_inst_7_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_15),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_7.READ_MODE = 1'b1;
defparam promx9_inst_7.BIT_WIDTH = 9;
defparam promx9_inst_7.RESET_MODE = "SYNC";
defparam promx9_inst_7.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_06 = 288'h4DA6D369B4DA6D369B4DA6D36DBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E9B4DA6D369B;
defparam promx9_inst_7.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_0F = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B6F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF9C;
defparam promx9_inst_7.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF7FBFBFDFEFFBFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_18 = 288'hFFFFFFE7D5DA6D369B4DA6D369B4DA6D369B4DA6D369BDE77FFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_20 = 288'hAF57ABD5EAF57ABD5EAF57ABD3E9F4FA3D1E7F379BCBE5F2F9BCFE8F4FA7D5EBF67F7FDF;
defparam promx9_inst_7.INIT_RAM_21 = 288'hAF57ABD5EAF57ABC9D6DA6D369B4DA6D369B4DA6D369B4DA6D369B5DC7ABD5EAF57ABD5E;
defparam promx9_inst_7.INIT_RAM_22 = 288'hFFE7EBF5EAF57ABD5EAF57ABD5EAF57ABD5EAF57ABD5EAF57ABD5EAF57ABD5EAF57ABD5E;
defparam promx9_inst_7.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_28 = 288'hBE7F53B3EDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_29 = 288'h7E3F1F8FC7E3F1F8FC7E3F1F8FC7E3F1F8DB4DA6CB67B2D9ECF67B3D9ECF67B2D9ED371C;
defparam promx9_inst_7.INIT_RAM_2A = 288'h7E3F1F8FC7E3F1F8FC7E3F1F8DB5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DAEDF8FC;
defparam promx9_inst_7.INIT_RAM_2B = 288'hFFFFFFFFFFF9F5F8FC7E3F1F8FC7E3F1F8FC7E3F1F8FC7E3F1F8FC7E3F1F8FC7E3F1F8FC;
defparam promx9_inst_7.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_31 = 288'h4DA6D36BB5DB6DB6FC8E670FB5FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_32 = 288'h4DA6D769B4DA6D369B4DA6D369B4DA6D369B5DAED369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_7.INIT_RAM_33 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_7.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFE7DF69B5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_7.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_3A = 288'h4DA6D369B4DA6D369B4DA6D369B4DAEE799C0EB7B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_7.INIT_RAM_3B = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6CF67B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_7.INIT_RAM_3C = 288'h3D9ECF67B3D9ECF67B3D9ECF67B3D9ECF67B3D9ECF67B3DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_7.INIT_RAM_3D = 288'hFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFC7A7B3D9ECF67B3D9ECF67B3D9ECF67B3D9ECF67B;
defparam promx9_inst_7.INIT_RAM_3E = 288'hEFE7F7F9FDFEFFFFDFEFFFFFFFFFFFFFBFFFEFF7FFFFFEFFFFFFFFFFF7F7FFFFFF7FBFFF;
defparam promx9_inst_7.INIT_RAM_3F = 288'hCFE7F3FBFFFF7F3FBFDFEFF3F9FFFF7F7FFFEFEFF7F9FCFE7FBFFFFFFFFFFBFDFEFFFFFF;

pROMX9 promx9_inst_8 (
    .DO({promx9_inst_8_dout_w[26:0],promx9_inst_8_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_17),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_8.READ_MODE = 1'b1;
defparam promx9_inst_8.BIT_WIDTH = 9;
defparam promx9_inst_8.RESET_MODE = "SYNC";
defparam promx9_inst_8.INIT_RAM_00 = 288'hFFFFEBD3EDFFFFFFFFFFFFFFFFFDFFFFFFFFFFF7FFFFFFFFFFFFBFCFE7F7FBFCFFFFFFBF;
defparam promx9_inst_8.INIT_RAM_01 = 288'hFFF7FFFFFFFFFFFFFFFFF7FBFFFFFFFFFFFFFFFFF3F9FDFFFFFFFFFFFFFBFDFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFDFFFFFFFFFFF7FFFFFEFFFFFFFFFFFFFBFDFEFE7F3F9FCFEFFFFFF;
defparam promx9_inst_8.INIT_RAM_03 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D367B5DDF0FB1EDFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_04 = 288'h4DA6D369B4DA6D369B4DA6DF7BCDE6F379BCDE6F379BCDE6F6F93C5DA6D369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_05 = 288'hAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE572B95CAE571369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_06 = 288'hFFDF9FDFFFFFFF3EDEFFFFFFFFFFFFFFFFFFFFFFEFF7CAE572B95CAE572B95CAE572B95C;
defparam promx9_inst_8.INIT_RAM_07 = 288'h6F2FA3DFFCFAF9BCBE6F2F77FDF5EF7FFFFFFFE7D7DFFBF47BFFFF8F67FFFFFFFCF93BDF;
defparam promx9_inst_8.INIT_RAM_08 = 288'h5F6FF3EDE5F2F97C9DFFE7D7ADE3E9F57CBEFFE7D3BFFDF9F5BCBE5F2FAFDFFFFDF97CDE;
defparam promx9_inst_8.INIT_RAM_09 = 288'hFFFFFFFFFFFB78FA9E5ED7BFFFFFFFFFFFFF5F77FFFFFFFAFBBFFFFFFFFFEDE5F274FABE;
defparam promx9_inst_8.INIT_RAM_0A = 288'h5F177BFFFDFA7BFFFFFFFFFFFFFFFC797DFFFFFFFFFFFBF3797CDE4F5FFFFFFFFFFDBCFE;
defparam promx9_inst_8.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFF5F67FFFFFFFC7ABDFF9F5FBFFFFFFFFDFD5ECF3797CBE;
defparam promx9_inst_8.INIT_RAM_0C = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6CF75C6F67FFFFF;
defparam promx9_inst_8.INIT_RAM_0D = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6EF9BFDFEFF7FBFDFEFF7FBFDFEFEBEBEBE36D369B;
defparam promx9_inst_8.INIT_RAM_0E = 288'h8F47A3D1E8F47A3D1E8F47A3D1E8F47A3D1E8F47A3D1E8F47A3D1E8F47A3D1E8F379369B;
defparam promx9_inst_8.INIT_RAM_0F = 288'hFF871F99FFFC7B7BFFFFFFEBD3CFFFFFFFFFFFFFFFFFFFFFFFFF5E9F47A3D1E8F47A3D1E;
defparam promx9_inst_8.INIT_RAM_10 = 288'hFF8F639DD2EF77BBFFBFFF43BFDFED727DDFAE5FFFFFFFFC7A79FF7F773FFFF0EAFBFFFF;
defparam promx9_inst_8.INIT_RAM_11 = 288'hEEEF577DDFEDFEBC1DFEFF7BADBEFD7BFBFDAE473BBDDDFD79F7FFBFC73381DFEFF63DFF;
defparam promx9_inst_8.INIT_RAM_12 = 288'hFFFFEB97CDFFFFFFFFFFBEFFABECE0773DFFFFFFFFFFFAE5FBFFFFFFD72BDFFFFFFFBE3D;
defparam promx9_inst_8.INIT_RAM_13 = 288'hAF077FBFDFEA6EFDFFCFBF3BFFFFFFFFFFFFFF875F9BFFFFFFFFFF2EC73FA3DBE277FFFF;
defparam promx9_inst_8.INIT_RAM_14 = 288'h4DEF37FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCE37BFFFFFF8F47BFF3E9F7FFFFFFFFF7A7D;
defparam promx9_inst_8.INIT_RAM_15 = 288'hEFB75F87B5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_16 = 288'hFFFFE389B4DA6D369B4DA6D369B4DA6D369B4DA6D77BFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_18 = 288'h6F7F7FFFFFFD71F71EFFE7F39BFFFFFFFEFCDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_19 = 288'hEFF7FFFFFEFA6E3DDFEFDFF39DFFFF7FBFDFDFFF5BDFF4F177FFFFFFC7AF9FFCFD73FFFF;
defparam promx9_inst_8.INIT_RAM_1A = 288'hFFFFFFFDFEFF7DF95FEFFFFFFDFEFF7F7F1CAF7FFBFDF8F7737FDFFFFFDF77FFFA76B9DF;
defparam promx9_inst_8.INIT_RAM_1B = 288'h6F6F7FFFFFFFFF7B5C9F7FFFFFFCFAEF7FFFEF874FBFFFFFFFFFFFFEBFBFFFFFF8F4BBFF;
defparam promx9_inst_8.INIT_RAM_1C = 288'hFFFFFBA9EFFF7FBFDFEFE717DFFFFBEE7DFFFFFFFFFFFFF976B83DFFFFFFFBFCE3FBBFDF;
defparam promx9_inst_8.INIT_RAM_1D = 288'h4DA6D369B4DB6EF8FEFFFFFFFFFFFFFFFFFFFFFFFFFFF6F077FFFFFFC7B39FFBFEF3BFFF;
defparam promx9_inst_8.INIT_RAM_1E = 288'hFFFFFFFFFFFEFDFD7C4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_1F = 288'hFFFFFFFFFFFFFCFA7B4DA6D369B4DA6D369B4DA6D369B4DA6D365DFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_21 = 288'hEFDF2FFFFBFBF3FFFFFFAEC3A9EFFEFFB95EFFFFFFFBD5EFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_22 = 288'hFFE7FBA7DFFFFFFFFFFFAEE7DFFFFEFF795EFFFFFFFFFFF9F4BBFFAFFF73FFFFFC7AF9FF;
defparam promx9_inst_8.INIT_RAM_23 = 288'hFFBFAB9FFFFFFFFFFFFFFFF78FEFFFFFFFFFFFFFFFFDD2EFFFFFFFBF6F33FFFFFFFF789E;
defparam promx9_inst_8.INIT_RAM_24 = 288'hEECFBFFFFBFC73FFFFFFFFF7A3D1EFFFFFFFEF8F7FFFFFFBFBFBDFFFFFFFFFF3EA7BFFFF;
defparam promx9_inst_8.INIT_RAM_25 = 288'hEF8753BFFFFFFFBA9EFFFFFFFFFFFA77BBFFFFFF57BFFFFFFFFFFFFF974FB5CCFFFFFFDF;
defparam promx9_inst_8.INIT_RAM_26 = 288'h4DA6D369B4DA6D369B4DA6D379C6F7FFFFFFFFFFFFFFFFFFFFFFFFAF777BFFFFFE7E79DF;
defparam promx9_inst_8.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFBEDE9D9ED369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFE7CDB4DA6D369B4DA6D369B4DA6D369B4DA6D371CEFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_2A = 288'hFFC7AF9FFFFFF4FBFFEFC733FFFDFA6DBC3DFFF7C3AFEFFFFFFE9ECE7FFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_2B = 288'hFFFFD7D9DFFFFE3DDDAF7FFFFFFFFF70BBFFFFF7FFAFEFFFFFFFFFFFB7BFBDFEF8F5BDFF;
defparam promx9_inst_8.INIT_RAM_2C = 288'h6F0F7FFFFFFE7D77DFFFFFFFFFFFFFFCBA7DFFFFFFFFFFFFFFFE9E9E7FFFFFFDFEF6BDFF;
defparam promx9_inst_8.INIT_RAM_2D = 288'h4F7FFFFFF1EB7BFFFFEFCF2FDFFFFFFF78DEFED7BFFFFFFDFFFFFFFFD7B79BFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_2E = 288'hFFF7EB93EFFCFAF9BFFFFFFBA9EFFFFFFFFFFFD7AB9BFFFAF87BFFFFFFFFFFFFF8F5BC5D;
defparam promx9_inst_8.INIT_RAM_2F = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369BAE47BBFFFFFFFFFFFFFFFFFFFFFCFF773FFF;
defparam promx9_inst_8.INIT_RAM_30 = 288'h9F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3EAED369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_31 = 288'h8F47A3D1E7F3FA3D5FEFFFFFFFFFFFFF7F7C4DA6D369B4DA6D369B4DA6D369B4DA6D765B;
defparam promx9_inst_8.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFDFDFCFE7F3FA3D1E8F47A3D1E8F47A3CFE8F47A3D1E8F47A3D1E;
defparam promx9_inst_8.INIT_RAM_33 = 288'hFFBFBFBFFFFC7AB9FFFFAFAB9FFFFF757DFFAF3F2BC1DDFFFCFA7EFFFFFFF7F6DF7FFFFF;
defparam promx9_inst_8.INIT_RAM_34 = 288'hEFFF5FDFFFFFFF3EFCEFFFFFE5D2EF7FFFFFFFCFB795EDFEFC7A9EFFFFFBF9FCFB7B39DF;
defparam promx9_inst_8.INIT_RAM_35 = 288'hFFFFFFFFF9F7777FFFFFFFDB75EFFFFFFFFFFFFFDBC1DEFFFFFFFFDFE7F3F1E4DF7FFFFF;
defparam promx9_inst_8.INIT_RAM_36 = 288'hFF8F5BDDFFEE7FFFFF7F176FFBFEFEF13BFFFFFFF7B1E5F0F7BFFFFFFFFFFFFDFA7B79BF;
defparam promx9_inst_8.INIT_RAM_37 = 288'hDFFF67DFFFFFFFFA5DFFFFEF8DEFFFFFFA9EFFFFFBF9FCFDFE797EFFCFBBBDFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_38 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B3DBF2BDFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_39 = 288'h4DA6D369BFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE71369B4DA6D369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_3A = 288'h4DAED76BB4DA6D369B4DA6D77BCBFFFFFFFFFFFFFFE3D4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_3B = 288'h5DDFFFFFFFFFFFFFFFFFFFFFFFFFF8F4F69B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_8.INIT_RAM_3C = 288'h4F176399FFFF7EB99FFFC7A79FFFFE7CF7FFFFB7BBBFF7F6773FFDCFFFDBDFDFFFFFFFFF;
defparam promx9_inst_8.INIT_RAM_3D = 288'h4DCFBFFFFFF9F4FDFFFFFFFFF1CBF7FFFF9FCE57FFFFFFFFFCFBDD7F4F87A1DFFFFE7C9E;
defparam promx9_inst_8.INIT_RAM_3E = 288'h5F470BBFFFFFFFFFFFCFEF33FFFFFFFFFA5DFFFFFFFFFFFFFEBDDDDFFFFFFFF7EA793C9E;
defparam promx9_inst_8.INIT_RAM_3F = 288'hFFFFFFFFFFF8F5BDFF3EB7BFFFFEF877F8FEAF07739FFFFFFF7B1EFFCEEFDFFFFFFFFFBF;

pROMX9 promx9_inst_9 (
    .DO({promx9_inst_9_dout_w[26:0],promx9_inst_9_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_19),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_9.READ_MODE = 1'b1;
defparam promx9_inst_9.BIT_WIDTH = 9;
defparam promx9_inst_9.RESET_MODE = "SYNC";
defparam promx9_inst_9.INIT_RAM_00 = 288'hFFFFFFFFFFF875BDFFFFFFDFD5CFFFFEBD7CFFFFC3A9EFFFFEBC7E4F2FAB8FEFFE7FBB9F;
defparam promx9_inst_9.INIT_RAM_01 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DAEEF97FFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_02 = 288'h4DA6D369B4DA6D369B9E67FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7DF89B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_03 = 288'h3DA6D369B4DA6D369B4DA6D369B4DA6D36BBDEEFFFFFFFFFFFFF1E6D9ED769B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_04 = 288'hEFFFFFFFFCE37BFFFFFFFFFFFFFFFFFFFFFFFFEFEB69B4DA6D369B4DA6D369B4DA6D367B;
defparam promx9_inst_9.INIT_RAM_05 = 288'hEFFFE7C9E4F27AB8DEFFFFDBB7CFFC7A79FFFFFFDB95FFFEFDF9FF2E9F7FFDDAF7FEBF9C;
defparam promx9_inst_9.INIT_RAM_06 = 288'h9F2793CBDAE1FBFFFFFFBFBBBFFFFFFFFFDD6F7FFFFFF7F573FFFFFFFFEFD9CDE077799C;
defparam promx9_inst_9.INIT_RAM_07 = 288'hFFFFE7D3CAE2F77FFFFFFFFFFFFEFF767DFFFFFFE3D9DFFFFFFFFFFFFFF3FBDBFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_08 = 288'hFFEFFB93EFFFFFFFFFFF975FDFF9F177BFFFFFDF9F7BC0EFF5B7DFFFFFF791EFFC787BFF;
defparam promx9_inst_9.INIT_RAM_09 = 288'hEFFFFFFFFFFFFFFFFFFF9F4BBFFFFFFF3EDBDFFFFFFFD7F7FC3A9EFFFFEFE9E4F27B7A9D;
defparam promx9_inst_9.INIT_RAM_0A = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B5DA6D761D;
defparam promx9_inst_9.INIT_RAM_0B = 288'h4DA6D369B4DA6D369B4DA6D369B6DB7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3A9B;
defparam promx9_inst_9.INIT_RAM_0C = 288'h5F2F97C7D9E26D369B4DA6D369B4DA6D369B4DA6D369B6DBFBFFFFFFFFFFFBFAE26D369B;
defparam promx9_inst_9.INIT_RAM_0D = 288'h5EFFF7F7CCFFFFFFFF4F077FFFFFFFFFFFFFFFFFFFFFFFFFFE3CBE5F2F97CBE5F2F97CBE;
defparam promx9_inst_9.INIT_RAM_0E = 288'h7F4FA3D5CDFFFF7F7FBFDFC7A1DFFFFF7F9C9F47A79FFFFFFF7A9EFFFFE397FEECFBFE3D;
defparam promx9_inst_9.INIT_RAM_0F = 288'h8F7FFFFFFDFDFEFF9F3EF77FFFFFFDFAB9FFFFFFFFE9E1EFFFFFFFDF8747BFFFFFFE7DBD;
defparam promx9_inst_9.INIT_RAM_10 = 288'h5F276F97EFFF7C3BFD7F67FFFFFFFFFFFFFFFF8F53DFFFFFFF7F5CEFFFFFFFFFFFFFBFDD;
defparam promx9_inst_9.INIT_RAM_11 = 288'hBFDFCFA1DFFF7C3ADEFFFFFFFFFFF8F43ABE3F572BDFFFFB7AF91E9F4F9F95EFFFFF383D;
defparam promx9_inst_9.INIT_RAM_12 = 288'h5DA6D36FC5EFFFFFFFFFFFFFFFFFFBFBBBFFFFFFFBF5B9F7FFFEDE2EF7FFA9EFFFFFBF7F;
defparam promx9_inst_9.INIT_RAM_13 = 288'hFFFFE3CDB4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_14 = 288'h1EA6D369B4DA6D369B4DA6D369B4DA6D369B4D877BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFBF4ECF1369B4DA6D369B4DA6D369B4DA6D369B4DF77FFFFFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_16 = 288'hBE6FFFEDEFEFFFFFDD7F7FFFFFFAF6F3BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_17 = 288'hFFFFE3DDDEFFFFFF9C9F7FFFFFFFFFFE3D3CFFFFFFEBE1EC7A79FFFFFFD7DDDFFFFFB8DE;
defparam promx9_inst_9.INIT_RAM_18 = 288'hFFFFFFE3D4F7FFFFFFFFFFFFFFFBF5F37FFFFFF7E797FFFFFFFF3EEEF7FFFFFFFD7B7B1E;
defparam promx9_inst_9.INIT_RAM_19 = 288'hFFFFF39FD3F2777ABEFFEFF78FEFFFFFFFDFCFFFFFFFFFFB7B79FFFFFFFFF9CBFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_1A = 288'hFFFFFFFFFFFFFE3DBCEFFFCFA5DFFFFF3FBFFF8F7B89E4F7747BFFFFAFB79FFFFFFF38BE;
defparam promx9_inst_9.INIT_RAM_1B = 288'h4DA6D369B4DA6D367B9DE7FFFFFFFFFFFFFFFFDFAF9FFFFFFFFFFC3EFFFFF9FFEDFFFA9E;
defparam promx9_inst_9.INIT_RAM_1C = 288'hFFFFFFFFFFFFFF3F7C4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_1D = 288'hFFFFFFFFF9F26D369B4DA6D369B4DA6D369B4DA6D369B4DD733FFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA75769B4DA6D369B4DA6D369B4DA6D369B4DB6F7FFF;
defparam promx9_inst_9.INIT_RAM_1F = 288'hEFFFD7C1DBE7FFFF7EAE7FFFE7DFE7FFFFFFDFE733FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_20 = 288'hFFFFD7DFDDFFFE7DDDDFFFFFE3D3EFFFFFFFFFFFF3EBCDFFFFFFDFDE2FA79FFFFFFF3F5C;
defparam promx9_inst_9.INIT_RAM_21 = 288'h6F7FFFFFFFFFFFFEBEFEFFFFFFFFFFFFFFFFEFD72FDFFFFFFF787DFFFFFFF9FDE67FFFFF;
defparam promx9_inst_9.INIT_RAM_22 = 288'hFFFFD3C1DFFFFF389DBFDFDBDFDEFEFFFB3EFFFFFFF7F4EFFFFFFFFFDF9F7DFFFFFFFE1D;
defparam promx9_inst_9.INIT_RAM_23 = 288'h2EB783A9EFFFFFFFFFFFFFEFF7CCFFFDFDBCFFFFE3D1EFF8F4BB7FBFCFAB99FFFC7AB9FF;
defparam promx9_inst_9.INIT_RAM_24 = 288'h4DA6D369B4DA6D369B4DA6D369B3DFF7FFFFFFFFFFFFFFFF7EF97FFFFFFFEBEFEFFFFFFF;
defparam promx9_inst_9.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFDD5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_26 = 288'h4D9ED3BFFFFFFFFFFFFFC71369B4DA6D369B4DA6D369B4DA6D369B4DA6E7DFFFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBA9B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_28 = 288'hFFFFFFF7CBFFFEBF3CDE7FFFFFF8E67FFF7F3DFFFFFFFEFEF2BFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_29 = 288'hFECFBFFFFFFFFFBFFD6F7FEFFFDCFFFFFEFEBE7FFFFFFFFFFFFEFB7F7FFFFFF4EFF279FF;
defparam promx9_inst_9.INIT_RAM_2A = 288'hFFFFFFE5D2EFFFFFFFFFFFFFF3E8DFFFFFFFFFFFFFFFFEFF75FDFFFFFFD3B5CFFFFFFFBF;
defparam promx9_inst_9.INIT_RAM_2B = 288'hFFEFD39FFFFFFEBD9DEFFFF791EFFFFFBFBDAF7FC7ABEFFFFFFF1E7E7FFFFFFFFFFDF75F;
defparam promx9_inst_9.INIT_RAM_2C = 288'hCE77FFFFFAF5F0789EFFFFFFFFFFFFFFBF9D9F7FEFF1BFFFFD7DDDFF8F5BDFFFFFFC7A3D;
defparam promx9_inst_9.INIT_RAM_2D = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DBF1FDFFFFFFFFFFFFFFFC3A3DFFFFFFF7F;
defparam promx9_inst_9.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7D5DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_2F = 288'h4DA6D369B4DA6E79FFFFFFFFFFFFFAF8F69B4DA6D369B4DA6D369B4DA6D369B4DA6FFBFF;
defparam promx9_inst_9.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7CFB4DA6D369B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_31 = 288'hAF571F9FFFFFFFFFFD7F7FF3F1CEEFFFFFFFDEAF7FFDFEE7F77FFFAF572BDFFFFFFFFFFF;
defparam promx9_inst_9.INIT_RAM_32 = 288'hEFFFFFFFF0EB7BFFDFBFE7F3EDEBE6FF7FDDBFFFFFF9F4DF7FFF9FBFE7F7FDC0EFFFFFFF;
defparam promx9_inst_9.INIT_RAM_33 = 288'hFFFFDFD5C9F7FFBF9C3EFFFFFFFFFFFFFFDF7E67FFFFFFFF7F3F9FCFFF4FBFFFFFFEFEBB;
defparam promx9_inst_9.INIT_RAM_34 = 288'hFFFFF3F5CCFFFD775FFFFFF7F9CBF7FF791EFFFFFFEDECE7FE7D7C8F77FBFFDAE7FFFFFF;
defparam promx9_inst_9.INIT_RAM_35 = 288'h6F77FFE5DCE7FFFFFFEF875B69EFFFFFFFBFBFDFF3FDC2EFFFBFDD2EFFD3D9CFF875BDFF;
defparam promx9_inst_9.INIT_RAM_36 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6FB9BFFFFFFFFFFFFFFEFF3C;
defparam promx9_inst_9.INIT_RAM_37 = 288'h4DA6DF79FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDE5DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_38 = 288'h4DA6D369B4DA6D369B4DA6D773EFFFFFFFFFFFE7DB69B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_9.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBE1D3DA6D369B;
defparam promx9_inst_9.INIT_RAM_3A = 288'hEEFFFFFFFEF87739FFFFFFFFE9E6F7FFBFFD3EFFFFFFF5F0F7FFFF9F0F4BA5DFE8777FFF;
defparam promx9_inst_9.INIT_RAM_3B = 288'hFFFFFBF3CBF7FFFFFF5F2F7FF9F2E974BA3DAE4FBBE1DBFFFFFFFF9E5FBFEFE2E974FBBC;
defparam promx9_inst_9.INIT_RAM_3C = 288'h5F7FFFFFFFFFFF7E5D2E9743BBD9F7FFFFFFFFFFFFFFFEEC7BFFFFFFCF8BA5D2EEF4FBFF;
defparam promx9_inst_9.INIT_RAM_3D = 288'hFF9F5FDFFFFFFFFE5D7F7FEB95EFFFFFBE1DAF7FFF93EFFFFFFFBFDE67FBE9E2E9747B9C;
defparam promx9_inst_9.INIT_RAM_3E = 288'hFFFFFFE9E2E9747BBC4EFFFFFFFFFCFA36DEFFFFFFF3E2E974BBBCFE7FFFF1E0E9777A7D;
defparam promx9_inst_9.INIT_RAM_3F = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6DF73EFFFFFFFFF;

pROMX9 promx9_inst_10 (
    .DO({promx9_inst_10_dout_w[26:0],promx9_inst_10_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_21),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_10.READ_MODE = 1'b1;
defparam promx9_inst_10.BIT_WIDTH = 9;
defparam promx9_inst_10.RESET_MODE = "SYNC";
defparam promx9_inst_10.INIT_RAM_00 = 288'h4DA6D369B4DA6CF6BEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1E6DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_01 = 288'h6DA6D369B4DA6D369B4DA6D369B4DA6D363DFFFFFFFFFFFFFF789B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_02 = 288'h0ECFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5E;
defparam promx9_inst_10.INIT_RAM_03 = 288'h2E974BA5D5F7FFFFFFFFCF97DFFFFFFFFF5E9F7FFFF1EAF7FFFFFFCFAFBFFFFFFD78BA1D;
defparam promx9_inst_10.INIT_RAM_04 = 288'h2E975FDFFFFFFFFE9ECFFFFFFFFAFCFBFF9F2E974BA5D2ECFBBEFEDFFFFFFFF5F67BFF1E;
defparam promx9_inst_10.INIT_RAM_05 = 288'h5E877FA5DEFFFFFFFFFFFFFFFBF3E877F8BEEFFFFFFFFFFFFFFFFF7F4FBFFFFFFCF8BA5D;
defparam promx9_inst_10.INIT_RAM_06 = 288'h6E8743B7FFFCFAFFFFFFFFFFF7E8F7FCFB9EFFFFFFF1EBFFFDBD9FFFFFFFFFF6F5FFFFDF;
defparam promx9_inst_10.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFF6F0743A5DCFFFFFFFFFFFFCFB5EFFFFFFF3E2E974BA5D4EFFFFFFF;
defparam promx9_inst_10.INIT_RAM_08 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6CF63D;
defparam promx9_inst_10.INIT_RAM_09 = 288'h4DA6D369B4DA6D369B4DA6D375CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1E6DA6D369B;
defparam promx9_inst_10.INIT_RAM_0A = 288'hFFFFFFFFFFEA6D369B4DA6D369B4DA6D369B4DA6D375CDFFFFFFFFFFFFDBCBB5DA6D369B;
defparam promx9_inst_10.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_10 = 288'h4DA6D36BBEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_11 = 288'h5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_12 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D36BBAF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFE;
defparam promx9_inst_10.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFCFB6D369B4DA6D369B4DA6D369B4DA6D36DC7F7FFFFFFFFFFEBD1C;
defparam promx9_inst_10.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_19 = 288'h4DA6D369B4DA6D369B2EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_1A = 288'hFFFFFFE9E5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_1B = 288'hFFFFFBFBC4DA6D369B4DA6D369B4DA6D369B4DA6D369B1EFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFEFEF5369B4DA6D369B4DA6D369B4DA6D369B1EFFFFFFF;
defparam promx9_inst_10.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFF5F7F77E3D9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_22 = 288'h4DA6D369B4DA6D369B4DA6D369B8E6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFE3D4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_24 = 288'hAE6FFFFFFFFFFFFE9D5DA6D369B4DA6D369B4DA6D369B4DA6D369BBE6FFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA79769B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFF7FEEBF83B9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_2B = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B3DC7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFBFBC4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_2D = 288'h4DA6D369B5DD7BFFFFFFFFFFF5E7E26D369B4DA6D369B4DA6D369B4DA6D369B7DC7BFFFF;
defparam promx9_inst_10.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7A389B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDE67379BFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_34 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DF77FFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_35 = 288'h4D9F7FFFFFFFFFFFFFFFFFFFFFFFFFFEFD3C4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_36 = 288'h4DA6D369B4DA6D369B3D8F7FFFFFFFFFFFFFCE26D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F389B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFC6CFBFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_3D = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DCF33FFFFFFFFFFFF;
defparam promx9_inst_10.INIT_RAM_3E = 288'h4DA6D369B4DDF3BFFFFFFFFFFFFFFFFFFFFFFFFFD7C9B5DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_10.INIT_RAM_3F = 288'h4DA6D369B4DA6D369B4DA6D369B4DB6FBFFFFFFFFFFFF8F1ED369B4DA6D369B4DA6D369B;

pROMX9 promx9_inst_11 (
    .DO({promx9_inst_11_dout_w[26:0],promx9_inst_11_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_23),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_11.READ_MODE = 1'b1;
defparam promx9_inst_11.BIT_WIDTH = 9;
defparam promx9_inst_11.RESET_MODE = "SYNC";
defparam promx9_inst_11.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFA9B;
defparam promx9_inst_11.INIT_RAM_01 = 288'hFFFFF7F7FBF5FAFD7FCFFFFFFFFFFFFFFFFFFFFFEFFDFFFFFFFFFFFFDFAFD7EBF5FB3DFF;
defparam promx9_inst_11.INIT_RAM_02 = 288'hFFE7EFD7EBFDFBBFFFFFFFFFF9FBFDFAFD7EBF5FBFFFFFFFFF3F7FEFFFFFFBFBFF7FFFFF;
defparam promx9_inst_11.INIT_RAM_03 = 288'hBF67FBFFFFFFFFFF7EBF5FAFD7FBFE7FFFFFFFFFFFFFFDFBF97D3EFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_04 = 288'hFFFFFFF9FCFFFFFFFFCFDFFFFFFFFFFFFFDFCFEFFFFFFFFDFB7FFFFFFFFFFFFBFDFAFD7E;
defparam promx9_inst_11.INIT_RAM_05 = 288'hFFFFFFF7ECFFFFFFFFFFF7EFD7FEFFFFFFBFCFFFFFFFFFFFFFFFFFBF1757B9FFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_06 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DB6E3DFF;
defparam promx9_inst_11.INIT_RAM_07 = 288'h4DA6D369B4DA6D369B4DAEEBDFFFFFFFFFFFFFFFFFFFFFFF7F389B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_08 = 288'hFFFFEBC9B4DA6D369B4DA6D369B4DA6D369B4D9EDBDFFFFFFFFFFFDFBF1369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_09 = 288'hBE5F3FBDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_0A = 288'hBE3FBFFFFFFFFE7D5CBE5F2F97C0EEFFFFFFFFFFFFFFFFFEFEF8DEFFFFFFFFFEFD72F97C;
defparam promx9_inst_11.INIT_RAM_0B = 288'hFFFFFFFFF5EE76F97CBE5F23DFFFFFFFFE5DBE673397CBE573BFFFFFFFE3D9D0EFFFFEFE;
defparam promx9_inst_11.INIT_RAM_0C = 288'hCE5F2F97CBE672BDFFFFFFFFFDDBE5F3397CBEF77FFFFFFFFFFF7EEED72795C0EE7FFFFF;
defparam promx9_inst_11.INIT_RAM_0D = 288'h5F7FFFFFFFFFFFFFFDEEE7FFFDF0EDF37FFFFFFFFFF5EDE27BFFFFFFE703BDFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_0E = 288'h4DAECFBFFFFFFFFFDDFEE7FFFFFFFFFD7B7C4EF7FFEBECE77FFFFFFFFFFFEBECE4F2799C;
defparam promx9_inst_11.INIT_RAM_0F = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_10 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6C7BFFFFFFFFFFFFFFFFFFFFFFAF9769B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFBEFC4DA6D369B4DA6D369B4DA6D369B4DA6F7BDFFFFFFFFFFFF875369B;
defparam promx9_inst_11.INIT_RAM_12 = 288'hEFBF2391C8E371B7DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_13 = 288'h5DAFBBEBE2D8F7FFFFFFFFE3CFC8E47238BB9E67FFFFFFFFFFFFFFFFEFCB61DFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_14 = 288'h6D9F77FFFFFFFFFFFFAE26DF71C8E1ECFDFFFFFFFFE3D7E470F69B7E3F33FFFFFFFEBD7C;
defparam promx9_inst_11.INIT_RAM_15 = 288'hFFFFFFFFFBE472391C7E1EDBDFFFFFFFFF9C7E3F0F6BB8E573FFFFFFFFFFE9D5DB6EB91C;
defparam promx9_inst_11.INIT_RAM_16 = 288'h3DCF278BB9E4FBFFFFFFFFFFF7C6E57FFF9F7E16E7DFFFFFFFFF3E6DEF7FFFFFFB6E799F;
defparam promx9_inst_11.INIT_RAM_17 = 288'h4DA6D369B4DA6FBBDFFFFFFFF5C7E57FFFFFFFFFDFD1CAE47BFE5D3DE7FFFFFFFFFF3D7C;
defparam promx9_inst_11.INIT_RAM_18 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_19 = 288'hFFCF9769B4DA6D369B4DA6D369B4DA6D369B4DA6DF7DFFFFFFFFFFFFFFFFFFFAFBF1369B;
defparam promx9_inst_11.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFE1D4DA6D369B4DA6D369B4DA6D369B4DAEDB95FFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_1B = 288'hEFFFFFFFFFF9F4FA7D3EEF1379FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_1C = 288'hFFFFFFF1E6DC72BD3E3DFF7FFFFFFFFF3E7D3E9F57D5C8DDFBFFFFFFFFFFFFFFFFFD77DD;
defparam promx9_inst_11.INIT_RAM_1D = 288'h4D8723C7D7E3727DFFFFFFFFFFF3DBF0BA9D2EBF03BFFFFFFFFF3E3F1F9373C2F1FB3FFF;
defparam promx9_inst_11.INIT_RAM_1E = 288'hFFD72395EFFFFFFFFF7F1F4FA7D1EA6D3DFFFFFFFFEFE3E875373C3F1F7FFFFFFFFFBF9C;
defparam promx9_inst_11.INIT_RAM_1F = 288'hFFFFE3CBB6DAF5BD9C4DF73BFFFFFFFFFE3D6E47BFF3E4DA6D7BFFFFFFFFF7F8E573FFFF;
defparam promx9_inst_11.INIT_RAM_20 = 288'h4DA6D369B4DA6D369B4DA6E79BFFFFFFFE1D6DC7BFFFFFFFFFFE9D6DF773EBE3DCFBFFFF;
defparam promx9_inst_11.INIT_RAM_21 = 288'h9E26D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_22 = 288'hFFFFFFFFFFFEFEF89B4DA6D369B4DA6D369B4DA6D369B4DA6CF6DEFFFFFFFFFFFFFFFF9F;
defparam promx9_inst_11.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF4DA6D369B4DA6D369B4DA6D369B4DA6D367D;
defparam promx9_inst_11.INIT_RAM_24 = 288'hFFFFE399CDFFFFFFFFFFFFFFFFFFFAF8F75EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_25 = 288'hDFFFFFFFFFFFFFFFFF6E9EF799F2DEF3FFFFFFFFFFFFFFFFFFFE5D6E57BFFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_26 = 288'hFFFFEFF1C7DFFFFFFF6E9EC3BFFFFFFFFFFF3DEF7BFFFBFCF2F9FFFFFFFFFFFFFFFDB79C;
defparam promx9_inst_11.INIT_RAM_27 = 288'hAE2EFFFFFFFFF5F73EFFFFFFFFFFFFFFFFFFCFBF03BFFFFFFFFFFFFFDFCF79CFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_28 = 288'h4DAF7FFFFFFFFDBC5B1EFFFFFBF8E3F27DFFFFFFFFEBE4DAFBFE3D4DA6C3BFFFFFFFFF9F;
defparam promx9_inst_11.INIT_RAM_29 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D777FFFFFFFE9E4DAFBFFFFFFFFFFFDF1E9EC3AFE;
defparam promx9_inst_11.INIT_RAM_2A = 288'hFFFFE7D9C5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_2B = 288'h4DA6D37BCEFFFFFFFFFFFFCBA9B4DA6D369B4DA6D369B4DA6D369B4DA6CF79CFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBE26D369B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_2D = 288'hFFFFFFFFFFFFFEF95CDFFFFFFFFFFF7EFF7FBF9F936BEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_2E = 288'hFFFFE793CBFFFFFFFFFFFFFFFFFDF975B83D6E5F3BFFFFFFFFFFDFBFDFEFE5D4DC7BFFFF;
defparam promx9_inst_11.INIT_RAM_2F = 288'hEFFFFFFFFFFFFEFEFCCE7FFFFFFDFC72F9BFFFFFFFFFF8E5733FFFDFDF1B7FFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_30 = 288'hFFFFFFFDFBE1EDFCFE8F77576FEFFFFFFFFFFFDFEFF7F9F4737BFFFFFFFFFFFFFF7D375C;
defparam promx9_inst_11.INIT_RAM_31 = 288'hCFE75B9FD6D8F7FFFFFFFFF7EDEBFFFFFFFF5F26D7DFFFFFFFFF5E3DA7BFF3C7DB6EF9FF;
defparam promx9_inst_11.INIT_RAM_32 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D36DEFFFFFFF3E3D9F7FFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_33 = 288'h8F57EBD5E7F17738BB4DA6D769B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_34 = 288'h4DA6D369B4DA6D371CAFFFFFFFFFFFFE3CDB4DA6D369B4DA6D369B4DA6D369B4DA6D36FC;
defparam promx9_inst_11.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4EA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_36 = 288'h3DB7BFFFFFFFFFFFFFFFFFFBAFCCFFFFFFFFFFE7FBB9DDED71363DFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFBAFCAF7FFFFFFFFFFFFFFFFFCF9771C5DD733FFFFFFFFFF7FCEE773B5C;
defparam promx9_inst_11.INIT_RAM_38 = 288'hFFFFDB71CCFFFFFFFFFFFFEFEFCEE7FFFFFFFFF71F97EFFFFFFFFF2EBEC3A9D3ECF137DF;
defparam promx9_inst_11.INIT_RAM_39 = 288'hDE4F1F9FFFFFFFFFFFDE1EEB95CBE47136DEFFFFFFFFFFF9773BBDCE2EEB9FFFFFFFFFFF;
defparam promx9_inst_11.INIT_RAM_3A = 288'hFFFFFFFFFFF8F4F6FC5DE73FFFFFFFFFFFDFFFFFFFFFFBF9EC7BFFFFFFFFFDF3D8F6FC9B;
defparam promx9_inst_11.INIT_RAM_3B = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D361DFFFFFFF9F3D8F7FFFF;
defparam promx9_inst_11.INIT_RAM_3C = 288'h4DA6D36BBDE077FBFDCE370F69B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_3D = 288'h4DA6D369B4DA6D369B4DA6D36BB4F7FFFFFFFFFFF7F5C4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_11.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAF3ED369B;
defparam promx9_inst_11.INIT_RAM_3F = 288'h7E3F1F8FC4D9F7FFFFFFFFFFFFFFFFFC7ABBBFFFFFFFFFFDFA78FC8E3F137BDFFFFFFFFF;

pROMX9 promx9_inst_12 (
    .DO({promx9_inst_12_dout_w[26:0],promx9_inst_12_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_25),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_12.READ_MODE = 1'b1;
defparam promx9_inst_12.BIT_WIDTH = 9;
defparam promx9_inst_12.RESET_MODE = "SYNC";
defparam promx9_inst_12.INIT_RAM_00 = 288'h7E2ECF79FFFFFFFFFFFFFFCBADB9F7FFFFFFFFFFFFFFFFFBF976DB3DC72BDFFFFFFFFF7F;
defparam promx9_inst_12.INIT_RAM_01 = 288'hFFFFFFFFFFFFFEB8FCAF7FFFFFFFFFFEFF1CCE7FFFFFFFF9F5373EFFFFFFFFFAF471B71C;
defparam promx9_inst_12.INIT_RAM_02 = 288'h4DFF53A7B4F5F137FFFFFFFFFFFFEA6DB8FC7E471367DFFFFFFFFFFFFF5F8FC7E2EDF9FF;
defparam promx9_inst_12.INIT_RAM_03 = 288'h5DFF7BFFFFFFFFFFFFEFFF4F6DB4DC73FFFFFFFFFFFFFFFFFFFFFFEFB6FBBDFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_04 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D377CFFFFFFFDF;
defparam promx9_inst_12.INIT_RAM_05 = 288'h4DA6D369B4DA6D369B3D9ECF67B3D9ECF67B3D9ECF67B3DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_06 = 288'hEFEF1369B4DA6D369B4DA6D369B4DA6D369BBE7FFFFFFFFFFFFE1D4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_08 = 288'hFFFFFFFDF5F2F97C7D6D877FFFFFFFFFFFFFFFFFD3C7BAF7FFFFFFFFF7DBCBE5F1F5F95C;
defparam promx9_inst_12.INIT_RAM_09 = 288'hDFE7136BB5E2ECF75EFFFFFFFFFFFFFDBA9B7F7FFFFFFFFFFFFFFFFFF7537FC4DBEE7DFF;
defparam promx9_inst_12.INIT_RAM_0A = 288'h4F5F137DFFFFFFFFFFFFFFFFADB8F7FFFFFFFFFFF7F7C8E7FFFFFFFFB78F6FEFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_0B = 288'hFFFFFFFFF7DEF738DBBFE70F7BFFFFFFFFFF3E9EFBABE5EA75363DFFFFFFFFFFFC797ABE;
defparam promx9_inst_12.INIT_RAM_0C = 288'hFFFFFFFFF7E6F3BFFFFFFFFFFFFCFBF137DC5DB6FFFFFFFFFFFFDFEFFFFFFFFFFC733BDF;
defparam promx9_inst_12.INIT_RAM_0D = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D371C;
defparam promx9_inst_12.INIT_RAM_0E = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6CB67B3D9ECF67B3D9ECF67B3D9ECF69B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_0F = 288'hFFFFFFFFFFF9F9769B4DA6D369B4DA6D369B4DA6D369B4DEFFFFFFFFFFFFF5E3DA6D369B;
defparam promx9_inst_12.INIT_RAM_10 = 288'hEFEFEF8BBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_11 = 288'h1EAEDFDFFFFFFFFFFFEFF7FBF9F9E6F7FFFFFFFFFFFFFFFFFE3C7B6F7FFFFFFFFFFFBFDF;
defparam promx9_inst_12.INIT_RAM_12 = 288'hFFFFFFFFFBF372B79FCF974F6DEFFFFFFFFFFFFFE7C7B5F7FFFFFFFFFFFFFFFDFAEE797F;
defparam promx9_inst_12.INIT_RAM_13 = 288'hFFF7FBFDFEF8F4F79FFFFFFFFFFFFFFCFA9B5F7FFFFFFFFFFFBFFD4DE7FFFFFFFB78F6FE;
defparam promx9_inst_12.INIT_RAM_14 = 288'hFFC72F9BFFFFFFFFFFCE471775CFFF74F75EFFFFFFFFF6E9EC3BDFEFEFE39DDEFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_15 = 288'h4DA6D36FCFFFFFFFFFAE5737FFFFFFFFFFFF5F2EE799FBE1EF7FFFFFFFFFEFE2EFFFFFFF;
defparam promx9_inst_12.INIT_RAM_16 = 288'h5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_17 = 288'hAE26D369B4DA6D369B4DA6D369B4DA6D369B4DCF0BA5D2E974BA5D2E974BA5D2E9743B7C;
defparam promx9_inst_12.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFDF9F89B4DA6D369B4DA6D369B4DA6D369B4D877FFFFFFFFFFFDF;
defparam promx9_inst_12.INIT_RAM_19 = 288'hFFFFFFFFFFFFFF387BDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_1A = 288'h2E9EFFBDF8F1ED7DFFFFFFFFFFFFFFFFFFBFCE4F3FFFFFFFFFFFFFFFFFE7CBB3EFFFFFFF;
defparam promx9_inst_12.INIT_RAM_1B = 288'hFF874F71EFFFFFFFFFBF373B9FFFFB75363DFFFFFFFFFFFFFEFE9B2EFFFFFFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_1C = 288'hEFFFFFFFFFFFFFFFFFFFA78F71EFFFFFFFFFFFFFE3C7B3F7FFFFFFFFFFFFEBE5DFF7BFFF;
defparam promx9_inst_12.INIT_RAM_1D = 288'h7E37BFFFFBFAEF39DFFFFFFFFFFEE2ECF63DFF974F6DEFFFFFFFFF9F26FBBFFFFF7EB97C;
defparam promx9_inst_12.INIT_RAM_1E = 288'h4DA6D369B4DA6D36FCFFFFFFFFFEEC733FFFFFFFFFFDFEE1ECFDFFDE9EEBDFFFFFFFFE5D;
defparam promx9_inst_12.INIT_RAM_1F = 288'hCFE7EBEDE1EDF1769B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_20 = 288'hFFFFFFFFF5F26D369B4DA6D369B4DA6D369B4DA6D369B4DCF33F9FCFE7F3F9FCFE7F3F9F;
defparam promx9_inst_12.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F389B4DA6D369B4DA6D369B4DA6D369B4DBF37FFF;
defparam promx9_inst_12.INIT_RAM_22 = 288'hFEFFFFFFFFFEFD7C9E4F27A787BAF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_23 = 288'hFFFFFFFDF9DAED7DFFBF9ECFBFFFFFFFFFBF4F2793C9DAE36FFFFFFFFFFBEBE4F2787ABB;
defparam promx9_inst_12.INIT_RAM_24 = 288'hAE3713B1E6F4F1B75EFFFFFFFFFCFBF379FFFFCF9779CFFFFFFFFFFFFFF3EDC0EFFFFFFF;
defparam promx9_inst_12.INIT_RAM_25 = 288'hFFF7F391CEFFFFFFFFFFC793C9E4F775367DFFFFFFFFFFFFFF3E7B1EFFFFFFFFFFFFFF7E;
defparam promx9_inst_12.INIT_RAM_26 = 288'hFFFFFFEFE5DDF1BCFE0E9EC3BDFFFFFFFFFF1E9ED373EFFAF8F65DFFFFFFFFFCFA6EF9FF;
defparam promx9_inst_12.INIT_RAM_27 = 288'h4DA6D369B4DA6D369B4DA6D36FCFFFFFFFFF1EAEEFFFFFFFFFFF7F9E2EEFFFF0E9EDFDFF;
defparam promx9_inst_12.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFB7B38BB4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_29 = 288'h4D9EDFDFFFFFFFFFFFEFBF1369B4DA6D369B4DA6D369B4DA6D369B4DA6F3FFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3C7B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_2B = 288'h6DB6DB69BBE7FFFFFFFFDFA78DB6DB6D767B6F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_2C = 288'hDEFFFFFFFFFFFFFF3E3DC72FFFFDFAEC3BFFFFFFFFF9F6DB6DB8FB5DA6F7FFFFFFFF3D1C;
defparam promx9_inst_12.INIT_RAM_2D = 288'hFFFFFFFFF3EB71B79C9E26F79BFFFFFFFFFFCFC72B9FFFFE79771CFFFFFFFFFFFFFF7F3C;
defparam promx9_inst_12.INIT_RAM_2E = 288'hEF9EE79DFFFFFC3ABBDFFFFFFFFFFFF5B6DB6DAECF7FDFFFFFFFFFFFFFFBE9BFEF7FFFFF;
defparam promx9_inst_12.INIT_RAM_2F = 288'h4E9ECFBFFFFFFFFFDFDE2F2395C4DB71BDFFFFFFFFFFF4F1EDF9FFFFC78F7DDFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_30 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D36FCFFFFFFFFF4F1EE7DFFFFFFFFEDE4DE73FFFF;
defparam promx9_inst_12.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3F5B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_32 = 288'h4DA6D369B4DA6FBBFFFFFFFFFFFFFFF4F6BB4DA6D369B4DA6D369B4DA6D369B4DA6C3BFF;
defparam promx9_inst_12.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBE9B4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_34 = 288'hFFFFF7F1C4DA6D369B7E7FFFFFFFFE7EB89B4DA6D367B4EFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_35 = 288'hFFFFF7F7C9E7FFFFFFFFFFFFE1D4DEF3FFFFEFBF37BDFFFFFFFFDF5DA6D369B4D9EEFDFF;
defparam promx9_inst_12.INIT_RAM_36 = 288'hDE77FFFFFFFFFFFFFFFF9F5365B3DB6E3DFFFFFFFFFFFCFC6E77FFFFEFDB6DCEFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_37 = 288'hFFFFFFFFFFFAEDF97FFFFFCFA9BBF7FFFFFFFF874F69B4DA6D373CFFFFFFFFFFFFFFFEFC;
defparam promx9_inst_12.INIT_RAM_38 = 288'h3DBFBFFFF6EA6C3BFFFFFFFFFFFFFE70F67B3DEF37FFFFFFFFFFFF7F26FBBFFFFE7CB79C;
defparam promx9_inst_12.INIT_RAM_39 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D36FCFFFFFFFFF7F1EDBDFFFFFFFFFBC;
defparam promx9_inst_12.INIT_RAM_3A = 288'h4DA6DB9BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FCE1ED36BB4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_3B = 288'h4DA6D369B4DA6D369B4DA6E395EFFFFFFFFFFFBF9769B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_12.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3DA6D369B;
defparam promx9_inst_12.INIT_RAM_3D = 288'hAF57FBFFFFFFFFBF7FAFD7EBF5EBFFFFFFFFFFFFEFD5EAFD7EBD5FDFFFFFFFFFFFFFFFFF;
defparam promx9_inst_12.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFF7FBFFFFFFFFFFFFFFF9FAFE7FFFFFFFDFB3FFFFFFFFFFFFAFD7EBF5E;
defparam promx9_inst_12.INIT_RAM_3F = 288'hFFFFFFF7FCFFFFFFFFFFFFFFFFFFFEFE7CDE5F57FBFFFFFFFFFFFFFFDFAFFFFFFFFEFF7E;

pROMX9 promx9_inst_13 (
    .DO({promx9_inst_13_dout_w[26:0],promx9_inst_13_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_27),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_13.READ_MODE = 1'b1;
defparam promx9_inst_13.BIT_WIDTH = 9;
defparam promx9_inst_13.RESET_MODE = "SYNC";
defparam promx9_inst_13.INIT_RAM_00 = 288'hFFFFEBF9FFFFFFFFFFFFD7EFDFFFFFFF7F5FFFFFFFFFFFFE7EBD5EAFD7ABD7FFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_01 = 288'hFFFFFFF9FAFF7FFFFFEFD7F3FFFFFFFFFFFFFFE7E3CBE7F67FFFFFFFFFFFFFFEFD7B3FFF;
defparam promx9_inst_13.INIT_RAM_02 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D373CFFFFFFFFFEFD7BBFFF;
defparam promx9_inst_13.INIT_RAM_03 = 288'h4DA6D369B4DA6D36DEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F4F1369B5DA6D369B;
defparam promx9_inst_13.INIT_RAM_04 = 288'h5DA6D369B4DA6D369B4DA6D369B4DA6D76BDFFFFFFFFFFFE7EB89B4DA6D369B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E;
defparam promx9_inst_13.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFBFEFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_0B = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D379CFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_0C = 288'h4DA6D369B4DA6D369B4DA6D37DDEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF975B69B;
defparam promx9_inst_13.INIT_RAM_0D = 288'hFFFFFFFDFAE26D369B4DA6D369B4DA6D369B4DA6D37DCEFFFFFFFFFFF7C3A9B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_14 = 288'hFFDFEB89B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D37FD;
defparam promx9_inst_13.INIT_RAM_15 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D375CCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFF2EA6D369B4DA6D369B4DA6D369B4DA6D36FBCFFFFFFFFFFFFDBCDB;
defparam promx9_inst_13.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_1C = 288'h4DA6CF63DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_1D = 288'hFFFFFFFFFFFFFCBA9B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_1E = 288'hFFFFF7F1C4DA6D369B4DA6D369B4DA6D369B4DA6D371CAF7FFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8F36D369B4DA6D369B4DA6D369B4DA6D369B7F7FFFFFF;
defparam promx9_inst_13.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_25 = 288'h4DA6D369B4DA6CF6BEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFEFEBB4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_27 = 288'hAE7FFFFFFFFFFFFE1D4DA6D369B4DA6D369B4DA6D369B4DA6D36DB7F7FFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFDF1369B4DA6D369B4DA6D369B4DA6D769B;
defparam promx9_inst_13.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_2E = 288'h4DA6D369B4DA6D369B4DA6D371EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7C4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_30 = 288'h4DA6D369B4DD7BFFFFFFFFFFF5E5DA6D369B4DA6D369B4DA6D369B4DA6D369B5F7FFFFFF;
defparam promx9_inst_13.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F5369B4DA6D369B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_32 = 288'hFFFFFFFFFFFF7F7FFFFFFFFFFDFDFEFF7FBFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_33 = 288'hFFF7FBFDFEFF7FBFDFFFFFFFFFFEFF7FFFFFFFF7FBFFFFFF7F7FDFFFF7F7FDFFFFFFFFBF;
defparam promx9_inst_13.INIT_RAM_34 = 288'hFFFFFFFDFFFFFFFFDFEFFFFFFFFFFFFFFFFFFFF7FBFDFEFF7FBFFFFFF7FBFDFEFF7FBFFF;
defparam promx9_inst_13.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F5FCFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_37 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D775EFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_38 = 288'h3EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7E3DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_39 = 288'h4DA6D369B4DA6D36BB3D977FFFFFFFFFFFFFBE26D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF9769B4DA6D369B;
defparam promx9_inst_13.INIT_RAM_3B = 288'hDFFFF7E9DBFFFFFFFFFFCF8FB3EFFFFFFF3E3F1F53C9E4F67BFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_13.INIT_RAM_3C = 288'h5F2F97DDFFFC797CBE4F2793AFEFFFFFFFFF9F2FB7FFFEFB7A3DFFFFE7D3CFEFFEFD3ADE;
defparam promx9_inst_13.INIT_RAM_3D = 288'hFFFFFFFFFFFFFF7E9DCFFFFFF3E4EEFFFFFFFFFFFFFFFCFAF97CBE5F2F97DFFEFB797CBE;
defparam promx9_inst_13.INIT_RAM_3E = 288'h6F67FFFFFFFFFFBF3E6F379BCDE9F7FFFFFFFFEFDBCFEFFFFFFFFFFFE7D3C1D1EBFBBFFF;
defparam promx9_inst_13.INIT_RAM_3F = 288'h6F67FFFBF7F5FBFFFFDFB7A7DFFDFB79BCDE6F37ABDFFFFE7DBDDFFFFFFFFFFFFFFFFF1E;

pROMX9 promx9_inst_14 (
    .DO({promx9_inst_14_dout_w[26:0],promx9_inst_14_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_29),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_14.READ_MODE = 1'b1;
defparam promx9_inst_14.BIT_WIDTH = 9;
defparam promx9_inst_14.RESET_MODE = "SYNC";
defparam promx9_inst_14.INIT_RAM_00 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6DF79FFFFFFFFFFFFFFFFEBD9F7FFFFBF;
defparam promx9_inst_14.INIT_RAM_01 = 288'h4DA6D369B1EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7E3DA6D369B4DA6D369B;
defparam promx9_inst_14.INIT_RAM_02 = 288'h4DA6D369B4DA6D369B4DA6D369B4DC73BFFFFFFFFFFFF5F1ED369B4DA6D369B4DA6D369B;
defparam promx9_inst_14.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE389B;
defparam promx9_inst_14.INIT_RAM_04 = 288'hFFE7DF6BC7F7FEBC7B4EFFFFFFFFFFF0B7BDFFFFFFE7D2D9ECF65B5DB77FFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_05 = 288'hDFC70F65B2D96D375EFFEF0F67B3D9ECB75CEFFFFFFFF1E2EE7DFFDFD72B9FFFFD79377C;
defparam promx9_inst_14.INIT_RAM_06 = 288'h3DB6E3DFFFFFFFFFFFFFFFE7C7B5F7FFFE3C1DB7BFFFFFFFFFFFFF6F16CB67B2D96CF79F;
defparam promx9_inst_14.INIT_RAM_07 = 288'hFFFFFFF3B2DA77FFFFFFFFEFF5C3D9ECF65BAE7FFFFFFFFB78F69BEFFFFFFFFFF9F5369B;
defparam promx9_inst_14.INIT_RAM_08 = 288'hBE77FFF5E4D9F7FF1E4DFF3FFFF8F16F7BFF9F16CF67B3D96FFBFFFFA78B77FFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_09 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6F39BFFFFFFFFFFFFFFFBE9B;
defparam promx9_inst_14.INIT_RAM_0A = 288'h4DA6D369B4DA6D369B1EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDF4DA6D369B;
defparam promx9_inst_14.INIT_RAM_0B = 288'hFFFFD3A7B5DA6D369B4DA6D369B4DA6D369B5DAEDBDFFFFFFFFFFFCFC71369B4DA6D369B;
defparam promx9_inst_14.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_0D = 288'hFFF7D791BEFFFF3F1B9E67F3EFC1EFFFFFFFFFEF0F6BBCFFFFFF5EDE777BB9C4D9F7FFFF;
defparam promx9_inst_14.INIT_RAM_0E = 288'h5DDF2BB7EFF8F339BCDE57136FEFFBFAF97C5DAEEF9BCEFFFFFFFF7F26DFDFFEFF7577FF;
defparam promx9_inst_14.INIT_RAM_0F = 288'hEFEF4F65D4F471B7BFFFFFFFFFFFFFFEFEFC1EFFFFEFE3D9F7FFFFFFFFFFFFFBFE7338DC;
defparam promx9_inst_14.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFF3C3DC73FFFFFFFFDBC9B7DE7338DC5DFFFFFFFFFB79367B4F7FFFFFF;
defparam promx9_inst_14.INIT_RAM_11 = 288'hFFFFFFF3CAE67FFF9F8E773FFBFAE2EFBFFF8F1EFFBFFDFD72F97CBE2EF7BDFFFBF9769E;
defparam promx9_inst_14.INIT_RAM_12 = 288'h5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6C3BFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_13 = 288'h4DA6D369B4DA6D369B4DA6D369B2EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_14 = 288'hFFFFFFFFFFFFFF3EDB4DA6D369B4DA6D369B4DA6D369B4DA6C3BDFFFFFFFFFFEFFF5369B;
defparam promx9_inst_14.INIT_RAM_15 = 288'h5D877FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_16 = 288'hFF8F4F7BFFFFFE78FCCFFFFFEBD8E6F2FD7CCE7FFFFFFFFDF1F6DB2EFFFFFDFAF57EBF3E;
defparam promx9_inst_14.INIT_RAM_17 = 288'hEFCFA7D9C7E37A7DDFFFDFA7D3E9F378F67DFFEFE7D1E7E3727D3EFFFFFFFFFCFA6D3BFF;
defparam promx9_inst_14.INIT_RAM_18 = 288'hBE77FFFFFEFF76397ECF974B6FEFFFFFFFFFFFFFF3F5CCE7FFFF7E4DEF3FFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_19 = 288'hFFCF9F7FDFFFFFFFFFFFFFFFEFC7E2EE3DFFFFFFDBC7B3ECFA7D9C4DE7FFFFFFFAF9B6FC;
defparam promx9_inst_14.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFD8E57BFFBFBE4F3FFFF2E9EDBDFF8F1EC7BFFFFCFA7D3E9F6F679BF;
defparam promx9_inst_14.INIT_RAM_1B = 288'hFFFFFFFFF5DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DAED7DFF;
defparam promx9_inst_14.INIT_RAM_1C = 288'hFFAF9769B4DA6D369B4DA6D369B4DA6D369B3EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFBC4DA6D369B4DA6D369B4DA6D369B4DA6EB97FFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_1E = 288'hFFFFFFFFF7E777BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_1F = 288'hEFB6C7BFFFFA79375EFFFFFB8BC9FFFFFFBF0EB6CBB9D8E7FFFFFFFFCF2B97C8E6FFFFFF;
defparam promx9_inst_14.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFE7D6E4FBFFFFFFFFFBFDFEFDFD37FDFFFFFFFFFAE2EFBFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_21 = 288'hFF9F5F81D5DC7BFFFFEFB793DFFEF974F65DFFFFFFFFFFFFFFBFBC7E7FFFFBF5DCF3BFFF;
defparam promx9_inst_14.INIT_RAM_22 = 288'hFF975B79FFFE7E393CFFFFFFFFFFFFFFFEBBDE3EFBBFFFFFFE3C9B6F7FFFE5D4DCFBFFFF;
defparam promx9_inst_14.INIT_RAM_23 = 288'h4DC72BDFFFFFFFFFFFFFFFFFE9E6E4FBFFDFEEAEFFFFF9F2EFBBFF8F1ECBBFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFDF4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_14.INIT_RAM_25 = 288'hFFFFFFFFFFFCFA389B4DA6D369B4DA6D369B4DA6D369B4F7FFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFE5DA6D369B4DA6D369B4DA6D369B4DA6D76DE;
defparam promx9_inst_14.INIT_RAM_27 = 288'h3DBFBFFFFFFC7A3D3E8E5F37FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_28 = 288'hFFFFFFFFFEFCF37BDFFFB7976BDFFFFD3A9C6F7FFFFFFCFC71777C5DF7FFFFFFFBF3787E;
defparam promx9_inst_14.INIT_RAM_29 = 288'h8E3EF3FFFFFFFFFFFFFFFFFFF1E4DB7BFFFFFFFFE3CDE6F2F937BDEFFFFFFFFDEA6EBFFF;
defparam promx9_inst_14.INIT_RAM_2A = 288'h3DA7BFFFFFF8F6395E5D8F7FFFFFFFFF7F5E6F570F63DFFFFFFFFFFFFFFFE1D4DF7FFFFF;
defparam promx9_inst_14.INIT_RAM_2B = 288'hFFF7E3D1E8F074F75FFFF7EB89BEFFFFFFFFFFFFFFE9B2EEF1799EFFFFEFF1C0EDFF3E7D;
defparam promx9_inst_14.INIT_RAM_2C = 288'h4DA6D369B4DDF3BFFFFFFFFFFFFFFFFFFF1E4DBFBFFFF1E9EF7FFFFFD71F99F7F1ECFDFF;
defparam promx9_inst_14.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFF5F3DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_14.INIT_RAM_2E = 288'h4DA6D37FCFFFFFFFFFFFEFEB89B5DA6D369B4DA6D369B4DA6D36BB6F7FFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9F9E26D369B4DA6D369B4DA6D369B;
defparam promx9_inst_14.INIT_RAM_30 = 288'hFFB73BBBF4DDF3FFFFCF9ECB65B4DCF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_31 = 288'h3E9EDBDFFFFFFFFFFFEFEF679DFFFD79B9FDFFFFEBE7B2EFFFFFFFFFD71367B3DE7FFFFF;
defparam promx9_inst_14.INIT_RAM_32 = 288'h3DD7BFFFFDE36EBDFFFFFFFFFFFFFFFFFF9F4DA77FFFFFFFFEF83B1D96D377CDFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_33 = 288'h4DF77BB9C4DFF7FFFFFF87239BFCE5733FFFFFFFDFD3C3D9ECB6BDFFFFFFFFFFFFFFFE7D;
defparam promx9_inst_14.INIT_RAM_34 = 288'h7F26D3DFFFFDFD363B1D9ECF6FEFFFFF385BCFFFFFFFFFFFFFBE7B3ECF8B67DFFFFFBE1D;
defparam promx9_inst_14.INIT_RAM_35 = 288'h4DA6D369B4DA6D369B3DAF7FFFFFFFFFFFFFFFFFFFF9F3DA77FFFF4EA6E3DFFFFB7938BE;
defparam promx9_inst_14.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1D4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_14.INIT_RAM_37 = 288'h4DA6D369B4DA6D36DCEFFFFFFFFFFEFEB87B5DA6D369B4DA6D369B4DA6D371CAF7FFFFFF;
defparam promx9_inst_14.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEA6D369B4DA6D369B;
defparam promx9_inst_14.INIT_RAM_39 = 288'h3DAF7FFFFDFA6FBBFF0EB6EBDFFEFE76B95C9E372BDFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_3A = 288'hBFFFFFFFF8F1ECFBFFFFFFFFFFFFF8F5B7BFFFEFE393CFFFFF7E9BFEFFFFFFFAF371771C;
defparam promx9_inst_14.INIT_RAM_3B = 288'hFFFFFFEDE5DB7BFFFF3EAF1FDFFFFFFFFFFFFFFFFFFDF6D8F7FFFFFFFFD7DBCDE6F6791C;
defparam promx9_inst_14.INIT_RAM_3C = 288'hEFFFFFF3E7DAED769B3DD73FFFFFFF76B9DF8F36E3DFFFFD7A78BB4DD70FBBFFFFFFFFFF;
defparam promx9_inst_14.INIT_RAM_3D = 288'hFFEFDF81D6F1EDFDFFFFEFFF99CCE571767DFFFFC7A7B8F7FFFFFFFFFFEFC9B4F77E79BD;
defparam promx9_inst_14.INIT_RAM_3E = 288'h4DA6D369B4DA6D369B4DA6D367B9E67FFFFFFFFFFFFFFFFFFFFFBF7E077FFFF7F2ECBBFF;
defparam promx9_inst_14.INIT_RAM_3F = 288'hDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3EFC4DA6D369B4DA6D369B4DA6D369B;

pROMX9 promx9_inst_15 (
    .DO({promx9_inst_15_dout_w[26:0],promx9_inst_15_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_31),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_15.READ_MODE = 1'b1;
defparam promx9_inst_15.BIT_WIDTH = 9;
defparam promx9_inst_15.RESET_MODE = "SYNC";
defparam promx9_inst_15.INIT_RAM_00 = 288'h4DA6D369B4DA6D369B4DA6D369B5F7FFFFFFFFCFA389B5DA6D369B4DA6D369B4DA6D377C;
defparam promx9_inst_15.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6F371369B;
defparam promx9_inst_15.INIT_RAM_02 = 288'h4EA6F385D5D877FFFFDF9EEB87DEEA6D3BFFFFC79FCFE3F26E3DFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_03 = 288'h9F4F8BADB9F7FFFFFFCF9EFFBFFFFFFFFFFFFFA79375EFFFFEB8BBEFFFFFEDCDEF7FFFFF;
defparam promx9_inst_15.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFF3E6DFF7FFFF8F1ECFDFFFFFFFFFFFFFFFFFFFF9E6F7BFFFFFFFF3F3E;
defparam promx9_inst_15.INIT_RAM_05 = 288'hEEAFAB91CAFFFFFF1E6DCEC7A3D7E473BFFFFFEF2387D2EAEC3BFFFFBF976FB2EBFB3FFF;
defparam promx9_inst_15.INIT_RAM_06 = 288'hAF37339FFFFFFC3B3C3E9EE3DFFFFF7E7D1E8F37A399CFFFFD7C5B4EFFE3CBDEFFFE3C7B;
defparam promx9_inst_15.INIT_RAM_07 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D36BB3EFFFFFFFFFFFFFFFFFFFFFFFDFBE673FFFF;
defparam promx9_inst_15.INIT_RAM_08 = 288'h4DA6D367DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7D7A9B4DA6D369B4DA6D369B;
defparam promx9_inst_15.INIT_RAM_09 = 288'h3EB71369B4DA6D369B4DA6D369B4DA6D369BAE3F9FD1E8F0F5769B4DA6D369B4DA6D369B;
defparam promx9_inst_15.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E8F479FCFE7F3F9FCFE7F379BCDE;
defparam promx9_inst_15.INIT_RAM_0B = 288'hBE6FFFFDFFE9ED7D7E8E5F3FFFFCF9EDB71C8E26F79BFFFFFFFFFFAFAED3BFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_0C = 288'hFFFFFFFFFFFFFE7C9B7F7FFFFFFFFA6F39DFFFFFFFFFFFFBF936DEFFFFFBA7BAF7FFFF3C;
defparam promx9_inst_15.INIT_RAM_0D = 288'hDFFFFBEBEAFFFFFFFFFFFFFFF9F7E4F3BFFFCF9EC7BFFFFFFFFFFFFFFFFFFFFDECF37FFF;
defparam promx9_inst_15.INIT_RAM_0E = 288'hBFFFDFC7B7E571F89B3EFFFFEDE5DFF3BFDFBE372FFFFFFDF1771C8DA6E39BFFFBF9779C;
defparam promx9_inst_15.INIT_RAM_0F = 288'hFEC73BFFFCFBF279FFFFFFE3CFCDEA6E7DFFFFFFFFFFFFFF7F38FCFFFFEBC5B0EFFCBB5C;
defparam promx9_inst_15.INIT_RAM_10 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D379CFFFFFFFFFFFFFFFFFFFFFFFFFDF;
defparam promx9_inst_15.INIT_RAM_11 = 288'h5DAED769B4DAEE399FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFAB89B5DA6D369B;
defparam promx9_inst_15.INIT_RAM_12 = 288'h7E3F1F8DB7E2ED369B4DA6D369B4DA6D369B4DA6D369B4DBF2393CAEB6D36BB5DAED76BB;
defparam promx9_inst_15.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDDAE4F2391C8E3F1F8FC;
defparam promx9_inst_15.INIT_RAM_14 = 288'h2EEFF7F3CAE67BFF9FAE26F7FDFAE36FFFFFAF9EDB71C8E3F1F95EFFFFFFFFFCFC703BFF;
defparam promx9_inst_15.INIT_RAM_15 = 288'h1EB6F3FFFFFFFFBF9FCFE7E7C9B4EFFFFFFFFFC72B99FFFFFF7F9FCFBF9B63DFFFFD3C7B;
defparam promx9_inst_15.INIT_RAM_16 = 288'hFFD7977BDDFF7E7C7B3EFFFFFFFFFFFFFFFFBE26E7DDFBF1EC3BFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_17 = 288'hBE77CBA7B8F7FD7C7B6E371F8BBBE77FFEFE5D8F7FFFF0EAEE7DFFEFCF176DB7E36CF6FE;
defparam promx9_inst_15.INIT_RAM_18 = 288'hFFFFFFFFF3EA6E7DDFBF3F1F7DFFFFFF7F7C6DA6EFDFFFFFFF7FBFDFE7F7A9BEFFFFBE5B;
defparam promx9_inst_15.INIT_RAM_19 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6E395EFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_1A = 288'h6DB6DB6DB6DB6DB6DB7E672FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF1369B;
defparam promx9_inst_15.INIT_RAM_1B = 288'h7E3F1F8FC7E3F1F8BB7E371369B4DA6D369B4DA6D369B4DA6D369B4DAEDF8FC7E36DB6DB;
defparam promx9_inst_15.INIT_RAM_1C = 288'hDFDF2F9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7C5DBF1F8FC;
defparam promx9_inst_15.INIT_RAM_1D = 288'hFFFFFBE9B6D8F43A9BBE6FFFF1E5DD6FFFFFCE1EF7FFF7F1EC7BBFDFCF9B85DFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_1E = 288'hFFFFFFFFF5F26EFFFFFFFFE3D5CAE56EB89B0EFFFFFFFFFFF6395EFFEFFFB5CAE4F1779C;
defparam promx9_inst_15.INIT_RAM_1F = 288'hDFD7A38FBFFFFEB8BB2EB7AB87B3EFFFFFFFFFFFFFFFF6F1EEB89DCE1EC3BFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_20 = 288'hBFFFFFF1B5E2FB789B6F7FCBABC6F6FF7E5D4DDFFFF5F6E673FFFF6EA6D7DFFEFB6F799E;
defparam promx9_inst_15.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFF9F3F238BD1E2EDF7FFFFFFFFE3D4DA6F3FFFFFF7CBBBDEEF76387B;
defparam promx9_inst_15.INIT_RAM_22 = 288'h0EB6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B3DBED7DDFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_23 = 288'h8F47A3D1E8F47A3D1E8F47A3D1E8F57BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9F;
defparam promx9_inst_15.INIT_RAM_24 = 288'h8F47A3D1E8F47A3D1E8F47A3D1E8F47A389B4DA6D369B4DA6D369B4DA6D369B4DCF1FD1E;
defparam promx9_inst_15.INIT_RAM_25 = 288'hFFFFFFFFFEFFF1B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E;
defparam promx9_inst_15.INIT_RAM_26 = 288'h5DAED36FBFFFFFFEBD7E371B69B1EFFFFE5D4D9F7FFFF1E9EE3DFF6F26D3DFFFFEFF391C;
defparam promx9_inst_15.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFF7F26DFDFFFFFFEFC9B5DAED769BCE7FFFFFFFFAF9771EFFF7FBABB;
defparam promx9_inst_15.INIT_RAM_28 = 288'hEFA6FFBFFFFF7FB87B8F7FE3D1B6E471371C9F7FFFFFFFFFFFFFFFDFF7576DC5DB71FDFF;
defparam promx9_inst_15.INIT_RAM_29 = 288'h5DAED367B5F7FFFEFE6E3F178DB9F7FFB8BB8F7FFFF3E6DEF3FF7F7E3F3FFFFBF16CBBFF;
defparam promx9_inst_15.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFEF8F576FC6D9EC7BFFFFFFFFF1E5D9EF7FFFFFF7FFA9B;
defparam promx9_inst_15.INIT_RAM_2B = 288'hFFEFDFC1D7E26D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B9E1F77FFF;
defparam promx9_inst_15.INIT_RAM_2C = 288'h4DC727DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7A7B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_15.INIT_RAM_2E = 288'hFFFFDBC3DFFFFFFFFFFFBF87BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_2F = 288'hFFF7DBC1D0E8743A3DFFFFFFFBF3EF77381DAF7FFFEFE0EDFBFFFF8F076FFFFAF0F67DFF;
defparam promx9_inst_15.INIT_RAM_30 = 288'hCE1773FFFFFFFFFFFFFFFFFFFFFBF8F6BDFFFFFFF7E1D0E8743A1D4EFFFFFFFFFDFC3B7F;
defparam promx9_inst_15.INIT_RAM_31 = 288'hEFFF5FDFFFFFF5BDFFFFFFE3DFD9F7FFFE9DEEE73789DDFFFFFFFFFFFFFFFFFFFCF83B9C;
defparam promx9_inst_15.INIT_RAM_32 = 288'hFFFFDBDDDFEFF7FBDD8F7FFFFDF2EE72F83DDFFFD3A1DBFFFFFFBF2E977FFBF1E8F7FFFF;
defparam promx9_inst_15.INIT_RAM_33 = 288'h4EF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD783B7CBE776BDFFFFFFFFFBF1EF77BFFF;
defparam promx9_inst_15.INIT_RAM_34 = 288'h9F4FA7D3E8F1F6F89B4DAED369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6DB75C;
defparam promx9_inst_15.INIT_RAM_35 = 288'h4DA6D369B4DAEC7B5EAFD7EBF5FAFD7EBF5FAFD7EBF5FAFCFA7D3E9F4FA7D3E9F4FA7D3E;
defparam promx9_inst_15.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFCBB4DA6D369B4DA6D369B;
defparam promx9_inst_15.INIT_RAM_37 = 288'hFFF7FFFFFFFFFFFFDFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_38 = 288'hFFFFFBFFFFFFFFBFDFEFF7FBFDFFFFFFFFFFFFE7E7D9FFFFFFFFDFEFFFFFFFFEFF7FFFFF;
defparam promx9_inst_15.INIT_RAM_39 = 288'hFFFFF7F3E9F77FFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFDFEFF7FBFDFEFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_3A = 288'hDFEFFFFFFFFEFFBFFFFFEFFBFFFFFFFFFFBFEFFFFFFFFCF4FA7FFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_3B = 288'hEFE7BFFFFFFFFFBFBFDFEFF7F9FEFFFFFFFFEFCF9FDBFFFFFF7FBFFFFFFFFFFEFEFFFFFF;
defparam promx9_inst_15.INIT_RAM_3C = 288'h4DAEF395FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF1E7F67FFFFFFFFFFFFFF;
defparam promx9_inst_15.INIT_RAM_3D = 288'h8E472391C8E47238FC4D9ED369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_15.INIT_RAM_3E = 288'h4DA6D369B4DA6D369B4DA6E39BCDE6F379BCDE6F379BCDE6F379BCCE472391C8E472391C;
defparam promx9_inst_15.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7C4DA6D369B;

pROM prom_inst_16 (
    .DO({prom_inst_16_dout_w[30:0],prom_inst_16_dout[9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_16.READ_MODE = 1'b1;
defparam prom_inst_16.BIT_WIDTH = 1;
defparam prom_inst_16.RESET_MODE = "SYNC";
defparam prom_inst_16.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_04 = 256'hFFFFFFFFFFFC000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_05 = 256'hFFFFE0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_06 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam prom_inst_16.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFF;
defparam prom_inst_16.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0E = 256'hFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0F = 256'hFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_10 = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_16.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFF;
defparam prom_inst_16.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_19 = 256'hFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1A = 256'hF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001F;
defparam prom_inst_16.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFF;
defparam prom_inst_16.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_23 = 256'hFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_24 = 256'hFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_25 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_16.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFF;
defparam prom_inst_16.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2D = 256'hFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2E = 256'hFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2F = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_16.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFF;
defparam prom_inst_16.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_37 = 256'hFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_38 = 256'hFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_16.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FF;
defparam prom_inst_16.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000003FFFFFFF;
defparam prom_inst_16.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000003FFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_17 (
    .DO({prom_inst_17_dout_w[30:0],prom_inst_17_dout[9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_17.READ_MODE = 1'b1;
defparam prom_inst_17.BIT_WIDTH = 1;
defparam prom_inst_17.RESET_MODE = "SYNC";
defparam prom_inst_17.INIT_RAM_00 = 256'hFFFFFFFFFFFFE0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_01 = 256'hDDEFFFFFFFFFFFFC0001FFF00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_02 = 256'hFFFFFFFFC0001FFFC00000003FFF7FFDC3BFDF97CF97F7BF070C0D93C9A37DBF;
defparam prom_inst_17.INIT_RAM_03 = 256'hFE0001FFFE00000001FFFFDBDFBBFDF7BCFBFF7FFDFEFBDDFBDFBFDBB9DEFFFF;
defparam prom_inst_17.INIT_RAM_04 = 256'hFFF00000000FFFBDFDFDBFEF7BDFFDFFDFDFEFBDDFBDFFBDBBBDEFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_05 = 256'h00007FFBDDDFDFFFFFBD7FDFFDFFFF7BEEFBDFDFDBBBFF7FFFFFFFFFFFE0000F;
defparam prom_inst_17.INIT_RAM_06 = 256'hBDDDFDDFF7FBDFFDFBDFFFF7BEFFDFFDDDDBBFF7FFFFFFFFFFFE0000FFFF8000;
defparam prom_inst_17.INIT_RAM_07 = 256'hFFFDDDBFBFBDFEFF7FEF7EFFDDDDDAEF7FFC0000000FF00007FFF800000003FF;
defparam prom_inst_17.INIT_RAM_08 = 256'hE7FBEFEFF7DEFBE4FDEDDDEEF7FFC00000007F00007FFFC00000001FFFEEFFDD;
defparam prom_inst_17.INIT_RAM_09 = 256'hFFBDFFFEEFFEDDD7EFFFFFFFF00007F00007FFFE00000001FFFEEFFDDFFFC9DF;
defparam prom_inst_17.INIT_RAM_0A = 256'hEEFEFDED76FBFFFFFF80003F80007FFFE00000000FFDEFDFFFFFBDDDDEFFFEFE;
defparam prom_inst_17.INIT_RAM_0B = 256'hF777BFFFFFFC0003F80003FFFE000000007FDEF5FEFFDBDDCDDFFDEFFFFBDF7D;
defparam prom_inst_17.INIT_RAM_0C = 256'hFFFFC0003F80003FFFE000000003FDF7FFEEFFDDFDEDFFDFFF7FBDF7EEFFEF5E;
defparam prom_inst_17.INIT_RAM_0D = 256'h01FC0001FFFF000000003FFF7BFEEEFFDEDEFF7DFFF7FBEF7EEF7EF9EE777BFF;
defparam prom_inst_17.INIT_RAM_0E = 256'h1FFFF000000001FEF7DFEEEFEDEDF6E7EEFF7FBEFFF6F7EF9EE773BFFFFFFE00;
defparam prom_inst_17.INIT_RAM_0F = 256'h0000001FFEFDFE7DFFDFDF7EFFEFF7FBEFFF7F7E7DFEFFF7FFFFFFF0001FC000;
defparam prom_inst_17.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFDFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FC0001FFFF00;
defparam prom_inst_17.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FE0000FFFF000000001;
defparam prom_inst_17.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FE0000FFFF000000000FFFFFFF;
defparam prom_inst_17.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FE0000FFFF000000000FFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFC0007F00007FFF0000000007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_15 = 256'hFFFFFFFFFFFFFC0007F00007FFE0000000007FFFFFF7FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_16 = 256'hFFFFFFC0007F00007FFE0000000003FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_17 = 256'h0003F80003FFE0000000003FFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_18 = 256'h003FFC0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_17.INIT_RAM_19 = 256'h000000003E7EF7F0FE7BF7BF03E03F0FF83F03EF7E0FFDF81FFFFFFFE0003F80;
defparam prom_inst_17.INIT_RAM_1A = 256'h01E7E77E07E73F39F03E03F07F03F03E77E07FDF81FFFFFFFE0001FC0003FFC0;
defparam prom_inst_17.INIT_RAM_1B = 256'hE63F73F39FFBFCFE73F3BFCFF33FE7FCFF9FFFFFFFF0001FC0001FF800000000;
defparam prom_inst_17.INIT_RAM_1C = 256'h39FFBFCFE7BF39FCFF93FF7FCFFDFFFFFFFF0001FC0001FF00000000001F7F37;
defparam prom_inst_17.INIT_RAM_1D = 256'hFE79F39FCFFD3FF7FCFFDFFFFFFFF0000FE0000FE00000000001F7FB7EF3F73F;
defparam prom_inst_17.INIT_RAM_1E = 256'hFCFFC3F07FCFC1FFFFFFFF8000FE0000FC00000000001F7F87FFBF61F39FF9FC;
defparam prom_inst_17.INIT_RAM_1F = 256'h07FEFC0FFFFFFFF8000FE00004000000000001F7FC3FFBF61F01FC1FCFE79FB9;
defparam prom_inst_17.INIT_RAM_20 = 256'hFFFFFFFF80007F00000000000000000F3F83FF9F29F01F81FCFE7DF81FEFFC3F;
defparam prom_inst_17.INIT_RAM_21 = 256'hFC0007F00000000000000000F3F83FF9F09F9DFF9FCFE7DF81FEFF83FF7FEFFC;
defparam prom_inst_17.INIT_RAM_22 = 256'h00003FFE000000000F3F93FF9F09FBCFFDFEFE7DF9DFEFF9BFF3FEFFCFFFFFFF;
defparam prom_inst_17.INIT_RAM_23 = 256'hF800000000F3F33F79F1DF9CFFDFEFF3DF9DFEFF9BFF3FEFFCFFFFFFFFC0007F;
defparam prom_inst_17.INIT_RAM_24 = 256'h000FBF3BF3BF9DF9CFF9FEFF39F9CFEFF3BFF3FE7FCFFFFFFFFC0003F80003FF;
defparam prom_inst_17.INIT_RAM_25 = 256'hBF03F9CF9EF80FE7F81F9CFE7F3BF03E07C0FFFFFFFFE0003F80003FFFC00000;
defparam prom_inst_17.INIT_RAM_26 = 256'hF9EFC0FE7FC3F9CFE7F39F03E07C0FFFFFFFFE0001F80003FFFE00000000FBF3;
defparam prom_inst_17.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FC0001FFFF00000000FBE7BF83F9C;
defparam prom_inst_17.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0001FC0001FFFF80000000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFF0000FE0000FFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2A = 256'hFFFFFFFFFF8000FE0000FFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2B = 256'hFFF8000FE0000FFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2C = 256'h7F0000FFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2D = 256'hFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_17.INIT_RAM_2E = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007F0000F;
defparam prom_inst_17.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007F0000FFFFF000;
defparam prom_inst_17.INIT_RAM_30 = 256'hE7E07CFC3FEF7F818180FB9CCEF8F07FFFFFFFFC0003F8000FFFFF0000001FFF;
defparam prom_inst_17.INIT_RAM_31 = 256'h99FEF7F81C1C0FB9CE6F8F07FFFFFFFFE0003F8000FFFFF0000001FE773981DF;
defparam prom_inst_17.INIT_RAM_32 = 256'hE7FDF3FBDCF278FF7FFFFFFFFE0003F8000FFFFF0000003FE733981DFE3E07CF;
defparam prom_inst_17.INIT_RAM_33 = 256'hBDCFA787F3FFFFFFFFE0001FC000FFFFF0000003FE73BBF9CFE3EE7C79DFE73F;
defparam prom_inst_17.INIT_RAM_34 = 256'h7F3FFFFFFFFF0001FC000FFFFF0000003FF739BFDCFE1EF7D7FDFE73FF7FCF3F;
defparam prom_inst_17.INIT_RAM_35 = 256'hFFFFF0000FC000FFFFF0000003FF7B9BFDCFE9EF7D7F9FF73FF7FCF3F9DEF879;
defparam prom_inst_17.INIT_RAM_36 = 256'h00FC000FFFFF0000007FF7BDBC1CFEDF03D3E1FF73FF7C0FBF9CEF879383FFFF;
defparam prom_inst_17.INIT_RAM_37 = 256'hFFFFE0000007FF7BDBC1EFECF039BC3FF7BFF7E0FBFDCE7879B83FFFFFFFFF00;
defparam prom_inst_17.INIT_RAM_38 = 256'h0000FFF39EBFCEFE4F339BCFFF3BFF3FEF9FDCE79793FBFFFFFFFFF8000FC000;
defparam prom_inst_17.INIT_RAM_39 = 256'h39E3FCEEE0F3381CFFF3BFF3FEF9FDCE73381FBFFFFFFFFF80007C001FFFFE00;
defparam prom_inst_17.INIT_RAM_3A = 256'h6E077B81CEFF3BFFBFEF9FDEE73381FBFFFFFE000000000001FFFFC000000FFF;
defparam prom_inst_17.INIT_RAM_3B = 256'hCCCFF93FFBE0F9C0E6733BDF9FFFFFE000000000003FFFF8000001FFFB9E3FCE;
defparam prom_inst_17.INIT_RAM_3C = 256'hFFBE07DC0F0F7BBCF9FFFFFFFFFC0003FFFFFFFF8000003FFF99F3E0E4EF73B9;
defparam prom_inst_17.INIT_RAM_3D = 256'hFFF9FFFFFFFFFFFFFFFFE0003FFFFFFFF0000007FFFC3F3C0F0CF33B9CE0FF83;
defparam prom_inst_17.INIT_RAM_3E = 256'hFFFFFFFFFFFFFE0003FFFFFFFC000000FFFFE3FBE0F9FFFFBBEF1FFE7FFFFFFF;
defparam prom_inst_17.INIT_RAM_3F = 256'hFFFFFFE000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_18 (
    .DO({prom_inst_18_dout_w[30:0],prom_inst_18_dout[10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_18.READ_MODE = 1'b1;
defparam prom_inst_18.BIT_WIDTH = 1;
defparam prom_inst_18.RESET_MODE = "SYNC";
defparam prom_inst_18.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_19 (
    .DO({prom_inst_19_dout_w[30:0],prom_inst_19_dout[10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_19.READ_MODE = 1'b1;
defparam prom_inst_19.BIT_WIDTH = 1;
defparam prom_inst_19.RESET_MODE = "SYNC";
defparam prom_inst_19.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_20 (
    .DO({prom_inst_20_dout_w[30:0],prom_inst_20_dout[11]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_20.READ_MODE = 1'b1;
defparam prom_inst_20.BIT_WIDTH = 1;
defparam prom_inst_20.RESET_MODE = "SYNC";
defparam prom_inst_20.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0DFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC093FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF801BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFA003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_04 = 256'hFFFFFFFFFFFA0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_05 = 256'hFFFFE000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_06 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_20.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFF;
defparam prom_inst_20.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFF40007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0E = 256'hFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0F = 256'hFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_20.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0002FFF;
defparam prom_inst_20.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00017FFFFFFFFF;
defparam prom_inst_20.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFF40001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_19 = 256'hFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1A = 256'hF00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001F;
defparam prom_inst_20.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0002FFFFFFFF;
defparam prom_inst_20.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFE80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_23 = 256'hFFFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_24 = 256'hFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_25 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_20.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFF;
defparam prom_inst_20.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0002FFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0002FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFD0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2D = 256'hFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2E = 256'hFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2F = 256'h00BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_20.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFF;
defparam prom_inst_20.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF40007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_37 = 256'hFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_38 = 256'hFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_39 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3A = 256'hFFF1CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_20.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000BFF;
defparam prom_inst_20.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFF00007FFFE1769A;
defparam prom_inst_20.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000010000400010001DFFFFFFF;
defparam prom_inst_20.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFA00000000000000000000015E7FFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3F = 256'hFBFB7DEF7E7F37B9EFFE0000000000000000000000007FFFFFFFFFFFFFFFFFFF;

pROM prom_inst_21 (
    .DO({prom_inst_21_dout_w[30:0],prom_inst_21_dout[11]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_21.READ_MODE = 1'b1;
defparam prom_inst_21.BIT_WIDTH = 1;
defparam prom_inst_21.RESET_MODE = "SYNC";
defparam prom_inst_21.INIT_RAM_00 = 256'hB4B79BFCFCFFF000000000400000030000000EFFFFFB7C7F7F9FFFCFCFF7FFFD;
defparam prom_inst_21.INIT_RAM_01 = 256'h8FCFFEFFFFFFFFFE0002003C00000013FFFBD3E05FF9F37DFD7F3DE9C2BF14FD;
defparam prom_inst_21.INIT_RAM_02 = 256'hFFFFFFFFE0000FFF00000000DFFF7B3C3D5FFFE7DFDDF79DE0C22BCDF306F9F3;
defparam prom_inst_21.INIT_RAM_03 = 256'hFC0001FFFE00000007FFFFBDE81FFDFC7F77DF7FE3624AAA30785F9B3AFC7FFF;
defparam prom_inst_21.INIT_RAM_04 = 256'hFFF00000003FFFD85EFFDFD63FE73EF3FFDFE79C8FBCFB197BDCE7FFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_05 = 256'h00007FF1B8EFBBFF773EBF9FFEFCFE7BFDF9BF819F1AAE7FFFFFFFFFFFF00007;
defparam prom_inst_21.INIT_RAM_06 = 256'h3FCEC7EFEBF1EBF9F7CFCF8B1E73EFC0BBFF7DF3FF800000007F00007FFF0000;
defparam prom_inst_21.INIT_RAM_07 = 256'hFFBB3EFF5F3FFEF97DE67DBE29FDB05FBFF80000000FE00007FFFC00000007FF;
defparam prom_inst_21.INIT_RAM_08 = 256'hEBF1CFCF9F9E73F546DBDA7D77FFE00000017F8000BFFFA00000003FFFCC4C78;
defparam prom_inst_21.INIT_RAM_09 = 256'h7EBDE7BEDF8EBED3673FFDFFF8000BF0000BFFFE000000017FFFECE1CFFDE8EF;
defparam prom_inst_21.INIT_RAM_0A = 256'hF6FEFBFEA6F9FFFFFF40007F00005FFFF00000000FFFEEADCDFD9EEDFB3F9F7D;
defparam prom_inst_21.INIT_RAM_0B = 256'h7F77DFFFFFFC0007F40001FFFD000000003FDF74FF6DC3DCD7EE7BE7E7F7BEBF;
defparam prom_inst_21.INIT_RAM_0C = 256'hFFFFA0001FC0001FFFE000000003F9F72FF7DE49CD3AF7EE7F7F3DFBCD7FCE5D;
defparam prom_inst_21.INIT_RAM_0D = 256'h02F80001FFFE800000001FCFB6FCCEFDDC4CEEFCFFF7FBCEFD777E7FEF7BF5FF;
defparam prom_inst_21.INIT_RAM_0E = 256'h0FFFE000000003FE2F4E055FC5DCEF1FCDFEBC5CFE166B271E57655FFFFFFD00;
defparam prom_inst_21.INIT_RAM_0F = 256'h0000002FF47EE968BE7C7F127DA7FFE5CF2607F477ECFFFFFFFFFFD0001F8000;
defparam prom_inst_21.INIT_RAM_10 = 256'hFF27CF873BFFECF6AFF27FBEBE72747647BEFF7FFFFFFFFE0001FE0001FFFE00;
defparam prom_inst_21.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FC0000FFFE000000000;
defparam prom_inst_21.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001FC00007FFF0000000017FFFFFF;
defparam prom_inst_21.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF4000FC0000FFFE8000000007FFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFF80007E80007FFF000000000FFFFFFEEFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_15 = 256'hFFFFFFFFFFFFFA000FF00003FFD0000000007FFFFFF8FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_16 = 256'hFFFFFF80003F00003FFF0000000007FFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_17 = 256'h0001F80005FFD0000000005FFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_18 = 256'h001FF80000000007E7877F4FE7FE3BF81E1BFFFF89E03D73F0FF8F81FFFFFFFC;
defparam prom_inst_21.INIT_RAM_19 = 256'h000000005E7EB3E4FE21E30F03F07FBBF01E03CB3E07F9F00FFFFFFFF0003F80;
defparam prom_inst_21.INIT_RAM_1A = 256'h02EBEB3C43EABE74F0BE13F6FF77E01D93C33F9F02FFFFFFFD0002FC0001FF80;
defparam prom_inst_21.INIT_RAM_1B = 256'hDFDF21F39FF7FDFF9DF23FC7EB3DFBFF7F8FFFFFFFF0002FE0001FF800000000;
defparam prom_inst_21.INIT_RAM_1C = 256'h3FFFDF8FEF3F1FFCFF23FE7FD7FDFFFFFFFF0002FE0000FE00000000003EBF47;
defparam prom_inst_21.INIT_RAM_1D = 256'h7DFBF5DFFFFF5EEFFCFBBFFFFFFFF8000FE0000FC80000000002EBE47EFFEB1E;
defparam prom_inst_21.INIT_RAM_1E = 256'hFE7FA1FE7FD7DBFFFFFFFF00017F00000800000000000F3F8BDF5E27E95FB3F9;
defparam prom_inst_21.INIT_RAM_1F = 256'h1BFE7A7FFFFFFFFC000FE00016800000000000E3FD7EFBF31F32FB7FE7FFFFE0;
defparam prom_inst_21.INIT_RAM_20 = 256'hFFFFFFFF00007F00000000000000000E9F93FF2F90F80F85FF7FFCF4CFDFF83F;
defparam prom_inst_21.INIT_RAM_21 = 256'hFE000BF00000000000000001FDF4BE7EF3CF3DF90FE7E7CFF8FF7FC3FEFFCF9A;
defparam prom_inst_21.INIT_RAM_22 = 256'h80007FFE000000001FFFA9F7BF0CF85F81FD7D3DFA6FE7FE1F03FCFC3FFFFFFF;
defparam prom_inst_21.INIT_RAM_23 = 256'h0600000001F9EB1FF2FDCFFA7FEFE7E1DFBFFDFF29FFBFE7FCFFFFFFFF80007E;
defparam prom_inst_21.INIT_RAM_24 = 256'h001F3F79EF1F9CF787D1FC7F06F18FDFF99F17D07E27FFFFFFFA0007F8000400;
defparam prom_inst_21.INIT_RAM_25 = 256'h5EE1F3DF4EFC0FD3FB1F7EFF7EFFF83D27C2FFFFFFFFC0001F40001FFF900000;
defparam prom_inst_21.INIT_RAM_26 = 256'hF8CFC1FF3F81F3D7C7FB2E03F0F807FFFFFFFC0003F80001FFFD00000001FBFF;
defparam prom_inst_21.INIT_RAM_27 = 256'hE7FD1FBCFFFE7DFFFFF7FFFFFFFFFFE0000FC0001FFFF80000001F1F33F03F9E;
defparam prom_inst_21.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0000FA0001FFFFC0000001F5EB1F97FDDF9F7BFF;
defparam prom_inst_21.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFE00007800017FFF40000001FFFFFFD7FFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2A = 256'hFFFFFFFFFF0001FE00007FFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2B = 256'hFFFC0007E00017FFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2C = 256'hFF0001FFFFE0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2D = 256'hFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_21.INIT_RAM_2E = 256'h0002FFFFFFFFFFFFFFFFFF7FEE7F818184F3DEAFFBEFFFFFFFFFF8000BF80017;
defparam prom_inst_21.INIT_RAM_2F = 256'h63D2DEFEBC37AF9BFDFFF00008FFF3CBFFFFF3FFFFFFFFE0003F0000FFFFF000;
defparam prom_inst_21.INIT_RAM_30 = 256'hE7F678FF3FC63F6638B373F99EFCEF3FFFFFFFFC0001F80007FFFF0000000FFF;
defparam prom_inst_21.INIT_RAM_31 = 256'h17FF6BFC0C5AF777B7179707FFFFFFFFC0001F40007FFFE0000001FCB231398F;
defparam prom_inst_21.INIT_RAM_32 = 256'h7EF9A3FBDC6779E9FFFFFFFFFC0000F4000FFFFF8000002FFEF11DCAFF7DBF87;
defparam prom_inst_21.INIT_RAM_33 = 256'hDBDF57CFF9FFFFFFFFF0003F8000FFFFF8000005FE7793B9DFFDCE7AB5DFDFBF;
defparam prom_inst_21.INIT_RAM_34 = 256'h363FFFFFFFFE8001FE000FFFFE0000007FF63D1FE9FEBDE7AB30FD61FF7C5F1F;
defparam prom_inst_21.INIT_RAM_35 = 256'hFFFFE8001FC0007FFFF0000001FFB923B98FE5F4B8FC8FE35FE7F971F0BC70BB;
defparam prom_inst_21.INIT_RAM_36 = 256'h007C0017FFFE0000003FE75D3A0E7EFD07FDE1FEB3FE3C1FDFC8CFC71F03FFFF;
defparam prom_inst_21.INIT_RAM_37 = 256'hFFFFC000000BFFFD97FEC7D9663ABB9FF7FFE7FAF7FBCE7271145FFFFFFFFE80;
defparam prom_inst_21.INIT_RAM_38 = 256'h0000FFEF1EDA4C546FC59BD1FFFDFF1DF71FCA6BE3B5B7FFFFFFFFF80007E000;
defparam prom_inst_21.INIT_RAM_39 = 256'h95CFF9C5E6733D1DD7F93FFBFE7CFAFE6B303F1FFFFFF607400034001FFFFA00;
defparam prom_inst_21.INIT_RAM_3A = 256'h468AF520D8FF41FF9C0F8E0EFA6304F5FFFFFF1F1400068007FFFFC000002FFE;
defparam prom_inst_21.INIT_RAM_3B = 256'hAF6FF3BFF1DAF8DAC0FF978FDFFFFFCFF8800078007FFFF0000000FFF28F5FA4;
defparam prom_inst_21.INIT_RAM_3C = 256'hFF5DCFA9DF9F715DF5FFFFFE7FEC0005FFFBFFFFC000002FFFD1F7B2745A2730;
defparam prom_inst_21.INIT_RAM_3D = 256'hE0F6E717EF9FFFFFFFFFE0003FFFFFFFE800000BFFF73FF9E62E67395A5AFFFD;
defparam prom_inst_21.INIT_RAM_3E = 256'hBEFDFFFFFFFFFE000400000001400001BFFF8DF1FF6DCFB71DEEEFFD9FFFE0FA;
defparam prom_inst_21.INIT_RAM_3F = 256'hFFFFFFE0002FFFBFFF000000EFFFFCBFBDE77FF7FDDFFCFFFBFF9E079C0FBE73;

pROM prom_inst_22 (
    .DO({prom_inst_22_dout_w[30:0],prom_inst_22_dout[12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_22.READ_MODE = 1'b1;
defparam prom_inst_22.BIT_WIDTH = 1;
defparam prom_inst_22.RESET_MODE = "SYNC";
defparam prom_inst_22.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA1FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80D7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE019FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFA007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_04 = 256'hFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_05 = 256'hFFFFD0013FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_06 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_22.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFF;
defparam prom_inst_22.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00017FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF40003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0E = 256'hFFFFFFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0F = 256'hFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_10 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_22.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFF;
defparam prom_inst_22.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00007FFFFFFFFF;
defparam prom_inst_22.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_19 = 256'hFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1A = 256'hF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0003F;
defparam prom_inst_22.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFF;
defparam prom_inst_22.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00017FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_23 = 256'hFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_24 = 256'hFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_25 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_22.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003FFFFFF;
defparam prom_inst_22.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFD00017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2D = 256'hFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2E = 256'hFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2F = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam prom_inst_22.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFF;
defparam prom_inst_22.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF40005FFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFC0002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_37 = 256'hFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_38 = 256'hFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3A = 256'hFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFF;
defparam prom_inst_22.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000018000C000018189;
defparam prom_inst_22.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFE0000C7FFFFFF;
defparam prom_inst_22.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFA0000000000000000000000C7FFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_3F = 256'h0C0D83F383FDFFDFFFFE0000000000000000000000079FFFFFFFFFFFFFFFFFFF;

pROM prom_inst_23 (
    .DO({prom_inst_23_dout_w[30:0],prom_inst_23_dout[12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_23.READ_MODE = 1'b1;
defparam prom_inst_23.BIT_WIDTH = 1;
defparam prom_inst_23.RESET_MODE = "SYNC";
defparam prom_inst_23.INIT_RAM_00 = 256'hB3079BF9FCFFE00000000040001FFD800000007FFF7FFF83BFFFC7FFF7FFBE06;
defparam prom_inst_23.INIT_RAM_01 = 256'hAFFFFF0000000000000000240000000BFFF3F7F7B7F9F97FFA3F7BF21D8CB73C;
defparam prom_inst_23.INIT_RAM_02 = 256'hFFFFFFFFE0000FFFC00000001FFF39FEBF3FCF3FF7A5F7FE3EFF57CD8B4DF9BB;
defparam prom_inst_23.INIT_RAM_03 = 256'hFE0000FFFA00000005FFF3BFEF9DFCEFBD717FF9FDFDF9F9FDCF9FBFFECF7FFF;
defparam prom_inst_23.INIT_RAM_04 = 256'hFFE800000007FF7BDEFD9FE7BFC7FFFFFFDFEF9CBF99FDDBFFF9E7FFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_05 = 256'h00007FF1E9EFCBFCF3FDFFCF79FFFE71DC79FFFBBBD0FEFFFFFFFFFFFFD0001F;
defparam prom_inst_23.INIT_RAM_06 = 256'hDCDEE79FD32DC3F0F1DFFF07FEE7B3E7F999D7FFFFFFFFFFFFFC00007FFFC000;
defparam prom_inst_23.INIT_RAM_07 = 256'hFDFBBCFEDF3FFC78BBEEBEBC4DBDD97FBFF80000000FE0000FFFFC00000007FF;
defparam prom_inst_23.INIT_RAM_08 = 256'hC1F9DFCF07FFFFE5E3FBF9E7F3FF800000003F8000BFFF800000001FFDCECE3A;
defparam prom_inst_23.INIT_RAM_09 = 256'h76BDE77C858D3EF2577FFDFFE8000FE8000FFFFE00000003FF9D7CE18FD3EDCF;
defparam prom_inst_23.INIT_RAM_0A = 256'hEF7EEBCD3EF7FFFFFE40003F80007FFFF000000007FDE76FFEFEFC1C5EBF9DFE;
defparam prom_inst_23.INIT_RAM_0B = 256'hD77F1FFFFFFE0005F00001FFFC000000003FFFFCFFFCC79CD6BF7FFFE7F9FEFB;
defparam prom_inst_23.INIT_RAM_0C = 256'hFFFFE0001F80001FFFE000000007FFE70FE6DDA9DDD4F7FEFEFFBFFBC4FFD79C;
defparam prom_inst_23.INIT_RAM_0D = 256'h01F80003FFFF000000003FCFF8FF5DDE9FCF6E7DE7E7FFDFBE77FF7BFD737BFF;
defparam prom_inst_23.INIT_RAM_0E = 256'h0FFFF800000000FFFFCF0EDDC5DCF477E77F387F7B00EE07BFDF3DFFFFFFFD00;
defparam prom_inst_23.INIT_RAM_0F = 256'h0000000FF87BE7E9FEEEEE3A7E27F39BEF283F7AFFE7F345FFFFFFF0000F8000;
defparam prom_inst_23.INIT_RAM_10 = 256'hFFB7FE77FBFFEEFF57ECFFF97E7A8B76B79F77393FFFFFFF0000FE0000FFFE80;
defparam prom_inst_23.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007C0001FFFE800000000;
defparam prom_inst_23.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8001FF0001FFFF800000000FFFFFFF;
defparam prom_inst_23.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007F0000FFFE000000000FFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFA0003F00003FFF000000000BFFFFFFEFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_15 = 256'hFFFFFFFFFFFFFC0003F00003FFF0000000007FFFFFFEFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_16 = 256'hFFFFFFE0003F80007FFF0000000003FFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_17 = 256'h0007F80003FFC0000000005FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_18 = 256'h007FFE0000000007E7CE7F8FE77F79F83F1BF4FF8BE03DE7D07FDF81FFFFFFFE;
defparam prom_inst_23.INIT_RAM_19 = 256'h000000003EBDEFED7FB5F3DFFDFFFF2BF7DFFDCFFDF3FAFFFFFFFFFFC0001F40;
defparam prom_inst_23.INIT_RAM_1A = 256'h01E7FA3D53F61E3CF71FCBF99F1BEDDFA3DF3F9FFBFFFFFFFE0003FC0001FFA0;
defparam prom_inst_23.INIT_RAM_1B = 256'hDA7E21FBFFF3F8FD15F0BEDDE03DC7FCFF8FFFFFFFF0003F80000FF000000000;
defparam prom_inst_23.INIT_RAM_1C = 256'h3CFF9F8FF7BF3DFF7FA7FF3FFFFCFFFFFFFE0001F80001FE80000000002EBF83;
defparam prom_inst_23.INIT_RAM_1D = 256'hFEF4F93FFFF03FF7FE7FCFFFFFFFF00007E0001FD00000000001E3F9BC61F21E;
defparam prom_inst_23.INIT_RAM_1E = 256'hFDFFB9FE3FE7D8FFFFFFFF8000FF00007B00000000001E7F9BCF1F77F33FB5FD;
defparam prom_inst_23.INIT_RAM_1F = 256'hE7FDFF8FFFFFFFF4000FC00007C00000000000E3F8FFFBE25F8CFFDFF7E79F2D;
defparam prom_inst_23.INIT_RAM_20 = 256'hFFFFFFFF8000FF00000000000000001F7FD7FFDF41F1DFFDFCFFFEFB0FF7FE7F;
defparam prom_inst_23.INIT_RAM_21 = 256'hFC0003F00000000000000000F7F27FFFF38F85F85FE7DF9F1DFCFF99F1FFC7E4;
defparam prom_inst_23.INIT_RAM_22 = 256'h00004003000000000F1F61FFCFEDF1AFF9FC7E39F81FC7F37FE3FE7F8FFFFFFF;
defparam prom_inst_23.INIT_RAM_23 = 256'h3800000000F5F3BE37F09F1DFFCFCFEFDF98FE7F99FEBFDFFE7FFFFFFFC0007F;
defparam prom_inst_23.INIT_RAM_24 = 256'h000F7FFBF1BF09F1DFF1FC7F2FF5BFDFEDBE97F1F82FFFFFFFFE0001F0000000;
defparam prom_inst_23.INIT_RAM_25 = 256'h3F75F38FBF7A5FEFFB0F5EFD7E33F89C2FC0FFFFFFFFC0003FC0001FFFE00000;
defparam prom_inst_23.INIT_RAM_26 = 256'hFEEFC1FE7FC1F78FF7F7DF03D07807FFFFFFFE0003FC0001FFFD00000000F9E7;
defparam prom_inst_23.INIT_RAM_27 = 256'hF7F87FFFFFFEFDF03F0FE07FFFFFFFF0003FE0000FFFF80000000FBE7FF85F3C;
defparam prom_inst_23.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE8002FA0000FFFFC0000001FBE7DF8FF1FFFCF81F;
defparam prom_inst_23.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFF0000FE0000FFFFA0000001FFFFFFEFFFFFFFFFFFFFFE7FF;
defparam prom_inst_23.INIT_RAM_2A = 256'hFFFFFFFFFF0000FD00007FFFC0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2B = 256'hFFFC000FC0000FFFFE0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2C = 256'hFF0001FFFFE0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2D = 256'hFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_23.INIT_RAM_2E = 256'h0001FFFFFFFFFFFFFFFFFD7FFFFFFFFFFBFFBDDEFDF07FFFFFFFF80007E00007;
defparam prom_inst_23.INIT_RAM_2F = 256'hEF153DFE3EC79F95FDEBF01C18FF1F9A5FAEF3FFFFFFFF80003F00007FFFF000;
defparam prom_inst_23.INIT_RAM_30 = 256'hE7F0787CBFC67F808380F11FACFCF0FFFFFFFFFC0003F00007FFFF0000000FE6;
defparam prom_inst_23.INIT_RAM_31 = 256'h82FE77FDF83F2F19EF078663FFFFFFFFC0007F00007FFFF0000002FEEFF303DF;
defparam prom_inst_23.INIT_RAM_32 = 256'h91C484FBCE6A7D767FFFFFFFFD0003F80007FFFF0000003FF2A713DEFF7EB787;
defparam prom_inst_23.INIT_RAM_33 = 256'h5CD61FDBF3FFFFFFFFF0003FA0007FFFF0000001FFEF33809FE5E13B7F1FCF7F;
defparam prom_inst_23.INIT_RAM_34 = 256'h7EDFFFFFFFFF0002F8000FFFFF0000001FF3713FABFF9C63CBBDFF7FFF3FCF7F;
defparam prom_inst_23.INIT_RAM_35 = 256'hFFFFE8000F8001FFFFF0000003FF79C3FCCFE3ED3BFF0FF71FEBE1F7F9EDF27B;
defparam prom_inst_23.INIT_RAM_36 = 256'h01F8000FFFFE0000003FE71E1C1C7C1E67E9E0FF71FE7E07BF9DEF87C707FFFF;
defparam prom_inst_23.INIT_RAM_37 = 256'h7FFFD000000BFE7FFB99C7EDE73DFE2FEBFFFFC3F3FABCF9393F7FFFFFFFFF00;
defparam prom_inst_23.INIT_RAM_38 = 256'h0001FFF79E9C2E4C07C3B7E5FEF3FF3C173FDFEFBB3BBBFFFFFFFFF400078000;
defparam prom_inst_23.INIT_RAM_39 = 256'h73D1FEEEE0ECBBEF7FE33FF1FCFBFDE6B1F3AFDFFFFFE7F8C00076000FFFFE00;
defparam prom_inst_23.INIT_RAM_3A = 256'h3496B5C1C47F1BFF1E0FCC5C1217A5F5FFFFFE207000024000FFFFE000001FFF;
defparam prom_inst_23.INIT_RAM_3B = 256'h5DE7FBBFF3D8FFBCE033101F3FFFFFE7FEC0003FFF7FFFFC000003FFF9BC3C2E;
defparam prom_inst_23.INIT_RAM_3C = 256'hFFBE2FAC1F06719AFBFFFFFEFFFE0003FFFFFFFEC000005FFF07F3CCE1F077D8;
defparam prom_inst_23.INIT_RAM_3D = 256'hDFEB7F7DDFFFFFFFFFFFC0001FFFFFFFB0000009FFF83F9FC7746739BC547F0F;
defparam prom_inst_23.INIT_RAM_3E = 256'hFFFFFFFFFFFFFF0001FFF8000E000003FFFFF3E7C0774E27FBF677FB9FFDDFFF;
defparam prom_inst_23.INIT_RAM_3F = 256'hFFFFFFF0000000C0010000001FFFFEBF3E0FACFB3BBE7BFFC7FFFFFFFFFF8FFF;

pROM prom_inst_24 (
    .DO({prom_inst_24_dout_w[30:0],prom_inst_24_dout[13]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_24.READ_MODE = 1'b1;
defparam prom_inst_24.BIT_WIDTH = 1;
defparam prom_inst_24.RESET_MODE = "SYNC";
defparam prom_inst_24.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC01FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8057FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFE004FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_04 = 256'hFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_05 = 256'hFFFFE000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_06 = 256'h0BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_24.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFF;
defparam prom_inst_24.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0002FFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0E = 256'hFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0F = 256'hFFFFFFA0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_10 = 256'h0002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_24.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFF;
defparam prom_inst_24.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_19 = 256'hFFFFFFFF40003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1A = 256'hFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0002F;
defparam prom_inst_24.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0001FFFFFFFF;
defparam prom_inst_24.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_23 = 256'hFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_24 = 256'hFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_25 = 256'h5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4000;
defparam prom_inst_24.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001FFFFFF;
defparam prom_inst_24.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80002FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2D = 256'hFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2E = 256'hFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2F = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE80;
defparam prom_inst_24.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFF;
defparam prom_inst_24.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_37 = 256'hFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_38 = 256'hFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_24.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FF;
defparam prom_inst_24.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000400001FF87;
defparam prom_inst_24.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000016FFFFFFF;
defparam prom_inst_24.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000038FFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFE000000000000000000000002FFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_25 (
    .DO({prom_inst_25_dout_w[30:0],prom_inst_25_dout[13]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_25.READ_MODE = 1'b1;
defparam prom_inst_25.BIT_WIDTH = 1;
defparam prom_inst_25.RESET_MODE = "SYNC";
defparam prom_inst_25.INIT_RAM_00 = 256'hFFFFF3BBBFFFC0000000004000200100000000FFFFFFFFFFFFFFFFFFCFFFFFFF;
defparam prom_inst_25.INIT_RAM_01 = 256'hBDDFFE00000000040001FFD00000000FFFFFD3EFBBFBF7BFFDBFFFFDFEF3DBDB;
defparam prom_inst_25.INIT_RAM_02 = 256'hFFFFFFFFE0001FFFE00000007FFFF93F39FFFF63CFF7F39ED8EB796DB5CDB9FF;
defparam prom_inst_25.INIT_RAM_03 = 256'hFC0000FFFE00000001FFFF93FFF9FCF7FF7FDFF9FEFF7FCDF99FF797F89FFFFF;
defparam prom_inst_25.INIT_RAM_04 = 256'hFFF80000000FFF3FFFFBFFCFB7E7BFF3FFFFF77FEF9EF979D7AEFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_05 = 256'h00007FFFE9FF9FFE77DFBBBFFDFCFF7DED7DFFFB9DFAFF7FFFFFFFFFFFC0001F;
defparam prom_inst_25.INIT_RAM_06 = 256'hDEDFFABFFF9BEBFFF7EFFFE7FDE78EFDF9DF1CE7FFBFFFFFFEFE00007FFF0000;
defparam prom_inst_25.INIT_RAM_07 = 256'hFF7B1EDFDFDEFDFF39F73DBDBCB9FFFF7FF800000017E0000FFFF800000001FF;
defparam prom_inst_25.INIT_RAM_08 = 256'hC7FDCFF773FFFFCEDFFBCF34FFFFC0000000FF0000FFFFE00000000FFFCCDDFF;
defparam prom_inst_25.INIT_RAM_09 = 256'h7979F7FD8E4E3DEAEFFFFC00080007F80007FFFE00000001FF9EFDDEEFF39FEF;
defparam prom_inst_25.INIT_RAM_0A = 256'hFE7EFBFF7FF3FFFFFFC0007F80007FFFE00000001FFFE77E1FFF1C2E8FFFBFFF;
defparam prom_inst_25.INIT_RAM_0B = 256'hF66FBFFFFFF80003F00003FFFE000000007F9F69FECFFFFFF9DFFDE7EFF3EE79;
defparam prom_inst_25.INIT_RAM_0C = 256'hFFFFC0003FC0001FFFF000000007FCFF5FCFDC39FE3EEF9EFFFF9CE7FDF7EF5E;
defparam prom_inst_25.INIT_RAM_0D = 256'h03FC0003FFFE000000007FCE71FE7FFCDCEE7EFEE7EFFFEFBFDF7E77E5FE7DFF;
defparam prom_inst_25.INIT_RAM_0E = 256'h3FFFF000000003FDE7FFF76FECE6F477E67FFFDCFFF777F73FFFFB5FFFFFFC00;
defparam prom_inst_25.INIT_RAM_0F = 256'h0000002FE1FBE0EABEEE6FE3FE37FB85E7F03731FDFF7B4FFFFFFFF0000FE000;
defparam prom_inst_25.INIT_RAM_10 = 256'hFFAFCE0FE9ECE7FBEFF7FFB83FF303FA0FBE77F9BFFFFFFE8000FC0001FFFE00;
defparam prom_inst_25.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FE0000FFFE000000000;
defparam prom_inst_25.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FD00007FFF000000000FFFFFFF;
defparam prom_inst_25.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80007E0000FFFF0000000007FFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFC0007E00007FFF000000000FFFFFFEFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_15 = 256'hFFFFFFFFFFFFFA0003E8000BFFE0000000007FFFFFE7FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_16 = 256'hFFFFFFC0003F00003FFD0000000007FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_17 = 256'h0003F80003FFE0000000007FFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_18 = 256'h001FFC0000000003FFFFFF3FFFBFFFF7FEE7FEFFF7FFFEFFEFFFFFFFFFFFFFFC;
defparam prom_inst_25.INIT_RAM_19 = 256'h000000001FFE77F4FFF3EF9F01E03EAFF81E03DF7C07FDF83FFFFFFFC0003FC0;
defparam prom_inst_25.INIT_RAM_1A = 256'h03EBFA7E43EB9EF9F7BECBE53F39ECFC73DE7FDFFDFFFFFFFF0001FC0001FFC0;
defparam prom_inst_25.INIT_RAM_1B = 256'hC63EA3EBAF81F13E09F57E13EC7E2BFDF85FFFFFFFF0000F80003FF400000000;
defparam prom_inst_25.INIT_RAM_1C = 256'h3EFF5FCFDFBF75FCFF93FEBFEFF8FFFFFFFF0000FC0001FF80000000003E3E73;
defparam prom_inst_25.INIT_RAM_1D = 256'hFD7DFB9FF7FABF07FCFC1FFFFFFFF0001FE0000FC00000000000F7F97E7DF61F;
defparam prom_inst_25.INIT_RAM_1E = 256'hFF7F93E07FFFA0FFFFFFFF00017E00010800000000001E3F73F7BE39F35FC7FD;
defparam prom_inst_25.INIT_RAM_1F = 256'hF3FC7BDFFFFFFFF00007E0000F000000000000F3F93FF3F0FF05F81FDFDFEF75;
defparam prom_inst_25.INIT_RAM_20 = 256'hFFFFFFFFC0007F00000000000000000F7FC7FFBF69FBCFFBFD7D78F59FC7FD5E;
defparam prom_inst_25.INIT_RAM_21 = 256'hF80007E00000000000000001FBFD3FFDFC1F39FB9FF7EFDF80FEFFD5FE7FE7FA;
defparam prom_inst_25.INIT_RAM_22 = 256'h00004002000000001F3FB3F7DF48F9FFF8FEFF7DF59FCFFA3FF7FEFFCFFFFFFF;
defparam prom_inst_25.INIT_RAM_23 = 256'hD800000001FFF91EF9F89F3CFF8FC7F7DF7CFC7F3BFF3FC7FCFFFFFFFFA0007F;
defparam prom_inst_25.INIT_RAM_24 = 256'h001F1E9BF3BF0CF9FFCCFE7E4CFF8FEFFB1F63ECFFE7FFFFFFFC0007F80007FF;
defparam prom_inst_25.INIT_RAM_25 = 256'h9F23F99FBEFD9FEFF43FD9FFFE5BE73FC79CFFFFFFFFE0003F80003FFFC00000;
defparam prom_inst_25.INIT_RAM_26 = 256'hFBC7C1FFFF85FFFFE7F3FF01F0FC0FFFFFFFFE0001FC0001FFFF00000001F1F3;
defparam prom_inst_25.INIT_RAM_27 = 256'hEFFDBF9CFE7F3BF03E07C0FFFFFFFFF0002FC0003FFFE00000001FBF7BFC3FB8;
defparam prom_inst_25.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE0001FE0001FFFFC0000001FBF7BFDBFBCF9EFC0F;
defparam prom_inst_25.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFF0001FE0001FFFF80000000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_2A = 256'hFFFFFFFFFF00017E0000FFFF80000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_2B = 256'hFFF8000FF00017FFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_2C = 256'hFF0000FFFFC0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_2D = 256'hFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_25.INIT_RAM_2E = 256'h0000FFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003E0000F;
defparam prom_inst_25.INIT_RAM_2F = 256'hBBDFDBFEFEF7FFF7FE67FFFFFB1F7FFDE78E0FFFFFFFFF80003F00007FFFE000;
defparam prom_inst_25.INIT_RAM_30 = 256'hE3D07CF87FCE7F8180C0F599DC7DE07FFFFFFFFE0007F80007FFFE0000003FF7;
defparam prom_inst_25.INIT_RAM_31 = 256'hCDFD73F20B9C1F3DDD77CEF3FFFFFFFFE0003FC0007FFFF0000001FE6371038F;
defparam prom_inst_25.INIT_RAM_32 = 256'h8D84C8F1DFF8FA707FFFFFFFFE0003FC0007FFFF0000003FF7F3383DFF7E47CF;
defparam prom_inst_25.INIT_RAM_33 = 256'h98E70FCFFFFFFFFFFFE0002FC0007FFFF0000003FFB73385BFF9E07D7A9FE63F;
defparam prom_inst_25.INIT_RAM_34 = 256'h7EBFFFFFFFFF0001FA0007FFFF0000005FEBB31F9FFE7CE3A3D8FEF7FEBF9F3F;
defparam prom_inst_25.INIT_RAM_35 = 256'hFFFFF8001FC000FFFFE0000003FF7BF1FCCFE0DA7A7E8FF7FFE7FCF9FBDEFC7C;
defparam prom_inst_25.INIT_RAM_36 = 256'h00FC0017FFFE0000007FF39D381CFE0F77F3E1FE3DFF3C0F3FDBCF83B785FFFF;
defparam prom_inst_25.INIT_RAM_37 = 256'hFFFFF000000FFFF9FBE0C7C4E83DBA1FF73FF7FF71F9FEF57B581FFFFFFFFF80;
defparam prom_inst_25.INIT_RAM_38 = 256'h00007FF37E1C7EDCD74FE3D7FE71FF7E07BF8EF703A9B3FFFFFFFFF8000FA000;
defparam prom_inst_25.INIT_RAM_39 = 256'hFFD9FDCC6A7759BCE7FBBFFBFCF9FDC67AB99F3FFFFFE7FF000074000FFFFC00;
defparam prom_inst_25.INIT_RAM_3A = 256'h466631DDBC7F13FF7FC7DFEE77331AFDFFFFFF3F8800060003FFFFA000000FFF;
defparam prom_inst_25.INIT_RAM_3B = 256'hAC67FA3FF9D8FEFDE87331AF9FFFFFE000000000009FFFFC000002FFF15E9FCE;
defparam prom_inst_25.INIT_RAM_3C = 256'hFFBC07CE0EE631BDFDFFFFFEFFFE0007FFFBFFFF8000003FFF71F1DE7ECE2BBF;
defparam prom_inst_25.INIT_RAM_3D = 256'hFFF57B55FFFFFFFFFFFFC0005FFFFFFFF800000BFFF9BF3E0FC76AF1BE5D7FD3;
defparam prom_inst_25.INIT_RAM_3E = 256'hFFFFFFFFFFFFFC0000000000080000017FFFA5F7FF71E737FFF78FFA3FF5FF7A;
defparam prom_inst_25.INIT_RAM_3F = 256'hFFFFFFE0003FFF7FFE0000000FFFFEFFFFFFBFFFFFFFF1FFE7FFFFFFFFFFDFFF;

pROM prom_inst_26 (
    .DO({prom_inst_26_dout_w[30:0],prom_inst_26_dout[14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_26.READ_MODE = 1'b1;
defparam prom_inst_26.BIT_WIDTH = 1;
defparam prom_inst_26.RESET_MODE = "SYNC";
defparam prom_inst_26.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0BFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF800BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_04 = 256'hFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_05 = 256'hFFFFC000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_06 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam prom_inst_26.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFF;
defparam prom_inst_26.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0E = 256'hFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0F = 256'hFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_10 = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_26.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFF;
defparam prom_inst_26.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_19 = 256'hFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_1A = 256'hFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001F;
defparam prom_inst_26.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFF;
defparam prom_inst_26.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_23 = 256'hFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_24 = 256'hFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_25 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_26.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFF;
defparam prom_inst_26.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_2D = 256'hFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_2E = 256'hFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_2F = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_26.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFF;
defparam prom_inst_26.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003FFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001FFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_37 = 256'hFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_38 = 256'hFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_39 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFF;
defparam prom_inst_26.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFE007F;
defparam prom_inst_26.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000DFFFFFFF;
defparam prom_inst_26.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000005FFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFE000000000000000000000001BFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_27 (
    .DO({prom_inst_27_dout_w[30:0],prom_inst_27_dout[14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_27.READ_MODE = 1'b1;
defparam prom_inst_27.BIT_WIDTH = 1;
defparam prom_inst_27.RESET_MODE = "SYNC";
defparam prom_inst_27.INIT_RAM_00 = 256'h1837DF7DDEFFFFFFFFFFFF80001FFE00000005FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_01 = 256'h9BEFFFFFFFFFFFF80003FFE800000017FFF7BFD83BFDF87CF87F7BE060C0D83C;
defparam prom_inst_27.INIT_RAM_02 = 256'hFFFFFFFFC0001FFF800000007FFFB93EBBBFDF2BFFAFFFFEDEEFBDAF97CB7F7B;
defparam prom_inst_27.INIT_RAM_03 = 256'hFC0000FFFD00000002FFF7FFEFDBFEFB7EFBDFB9FDFEF7DBFBFFD7FB7DFEFFFF;
defparam prom_inst_27.INIT_RAM_04 = 256'hFFE000000017FFFDDEFBDFDFFBE7BBF39FEFF7FEEFBFF9FFBBAFF7FFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_05 = 256'h0000BFFFDFEFFBFC73BEFFFF7DFCFEFFDFFDEFB9FDB8EEFFFFFFFFFFFFE0000F;
defparam prom_inst_27.INIT_RAM_06 = 256'hFEEEFDFFDF3DF3FBFFDFDFF7DEE7FEFBBFBDBCF7FFC0000001FF0000FFFF0000;
defparam prom_inst_27.INIT_RAM_07 = 256'hFD3ABFBF1FFEFFF079EFFD7E1FDDB7DF7FF80000001FE0000FFFFC00000003FF;
defparam prom_inst_27.INIT_RAM_08 = 256'hFBFFFFFF8BBF73FFE0CDDD3FFBFFE0000000FE00007FFFC00000003FFDFFCE0F;
defparam prom_inst_27.INIT_RAM_09 = 256'hFF7FE7FF7FCFDEDE7F7FFE00000003F00003FFFE00000001FF9EF4E2FFDBDDFB;
defparam prom_inst_27.INIT_RAM_0A = 256'hDFFDEDDEEF7FFFFFFF00007F80007FFFC000000007FBFE6FDEFE7BDE3F7F9EFF;
defparam prom_inst_27.INIT_RAM_0B = 256'hDFEFFFFFFFF80003F80007FFFF00000000FFFF7CFDCFE7BEF2EFFBFFE7FFDFFE;
defparam prom_inst_27.INIT_RAM_0C = 256'hFFFFE0001F80003FFFF000000007FFEF0FFDEDDFDEDFF7DE7EFFFEFFDFF7EFBF;
defparam prom_inst_27.INIT_RAM_0D = 256'h01F80003FFFE000000001FCFFCFFEDDCDFFFEF7DE7F7FDDFFF7EFEF5FEF77FFF;
defparam prom_inst_27.INIT_RAM_0E = 256'h1FFFE000000003FE6FCFF75DFDFFEFFFDF7F7FDEFBEFF7F7DF6FBFBFFFFFFE00;
defparam prom_inst_27.INIT_RAM_0F = 256'h0000001FE17CF1FA9E5EFFE37E3FFFC5FF30FFE1FFE773CFFFFFFFF0001FC000;
defparam prom_inst_27.INIT_RAM_10 = 256'hFF2FDF077FF5FDF76FF6FF7C1EFF06F707DFEFBDFFFFFFFF0000FE0000FFFF00;
defparam prom_inst_27.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8001FC0001FFFF000000000;
defparam prom_inst_27.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007E0000FFFE000000000FFFFFFF;
defparam prom_inst_27.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007F0000FFFE0000000007FFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFF8000FE0000FFFF0000000007FFFFFF5FFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_15 = 256'hFFFFFFFFFFFFFC0007F00007FFF0000000003FFFFFFBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_16 = 256'hFFFFFFE0003F80003FFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_17 = 256'h0003F00007FFC0000000003FFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_18 = 256'h003FFE0000000001FFFFFF9FFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_27.INIT_RAM_19 = 256'h000000001FFD6FEB7FF7FBDFFFFFFFDFF7FEFFFEBFF7FEFFFFFFFFFFE0001F80;
defparam prom_inst_27.INIT_RAM_1A = 256'h03F7C67F2FF73F7BF81F07E23F81E03F23E0FFDF81FFFFFFFE0003FC0001FF80;
defparam prom_inst_27.INIT_RAM_1B = 256'hE17E71F7DF01E03F23F03F03F37E17FDF85FFFFFFFF0001FC0001FF800000000;
defparam prom_inst_27.INIT_RAM_1C = 256'hBDFF9FDFE73F7BFDFF37FE7FDFF9FFFFFFFF0000FE0000FF00000000001E7E67;
defparam prom_inst_27.INIT_RAM_1D = 256'hFEFBF7DFCFF87FE3FFFF8FFFFFFFF8001FE0001FF00000000001E3F83C73E21F;
defparam prom_inst_27.INIT_RAM_1E = 256'hFEFFC7FF3FEFFCFFFFFFFF0000FC0000F200000000000F3FD3EF1F23F8CFFBFC;
defparam prom_inst_27.INIT_RAM_1F = 256'h03FCFC1FFFFFFFF80007F0000F800000000000F3F87FFBF29FB8FBBFCFEFDF21;
defparam prom_inst_27.INIT_RAM_20 = 256'hFFFFFFFFC000FF00000000000000001F7FC3FFBF45F80FC1FEFEF9F81FCFF83F;
defparam prom_inst_27.INIT_RAM_21 = 256'hF80007F00000000000000000F7F93FFBF6DF21FC5FEFF78FC1FC7FD3F07FCFC1;
defparam prom_inst_27.INIT_RAM_22 = 256'h80000003000000000FFF1BE7BF9DF1DFF9FC7F78FB8FE7F91FFFFC7FEFFFFFFF;
defparam prom_inst_27.INIT_RAM_23 = 256'hEC00000000FBF9BE3BF88FBFFF9FE7E7CFB8FE7F31FFFFE7FEFFFFFFFFC0007F;
defparam prom_inst_27.INIT_RAM_24 = 256'h000F3F39E4BF18FBEF84FE7F91FBDFEFF19F0BE0FC0FFFFFFFFE0003F00003FF;
defparam prom_inst_27.INIT_RAM_25 = 256'h1F91F1DF9EFC1FEFF1BFBCFEFF3BF03E0FE07FFFFFFFC0001F80003FFFA00000;
defparam prom_inst_27.INIT_RAM_26 = 256'hF9CFC0FEFF83F9CFFFF7BF03E07E07FFFFFFFE0003FC0001FFFE00000000F3E7;
defparam prom_inst_27.INIT_RAM_27 = 256'hFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFF0001F80001FFFF80000000F1F33FC7F3D;
defparam prom_inst_27.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0000FC0000FFFF00000000FFFFFFE7FFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFF8001FE0001FFFF80000001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2A = 256'hFFFFFFFFFF0000FC0001FFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2B = 256'hFFF00007E0000FFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2C = 256'h7F00007FFFE0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2D = 256'hFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_27.INIT_RAM_2E = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007F00007;
defparam prom_inst_27.INIT_RAM_2F = 256'h77B83DFF7F0FCFD3FEF7F8181C0FB9CCEFDF07FFFFFFFFC0003F80007FFFE000;
defparam prom_inst_27.INIT_RAM_30 = 256'hF3E0F8F81FE63F01C1C1F3FCC67DE03FFFFFFFFC0003F00007FFFF0000001FEF;
defparam prom_inst_27.INIT_RAM_31 = 256'hC1FE63FE7BCB3F9DCEE7CFF3FFFFFFFFC0001F80007FFFF0000003FEF27B839F;
defparam prom_inst_27.INIT_RAM_32 = 256'hF3F8F3F9DCE7FC7F7FFFFFFFFE0003FC0007FFFF0000003FEF7BBFB8FE3C6787;
defparam prom_inst_27.INIT_RAM_33 = 256'h99EF17B7F7FFFFFFFFF0001F80007FFFF0000001FF7B1BFFDFE3C778FD8FFF7F;
defparam prom_inst_27.INIT_RAM_34 = 256'h397FFFFFFFFE0000FC0007FFFF0000003FE7BB9F9CFEBE678798FF73FE7FDFBF;
defparam prom_inst_27.INIT_RAM_35 = 256'hFFFFF0001FE0007FFFF0000007FE3B99C5EFE5EE397F4FF73FF3C1FBFF8C797A;
defparam prom_inst_27.INIT_RAM_36 = 256'h00FE000FFFFE0000003FF3389C0EFE4F77DFD0FE7BFF3E1F1FFDEFC7B383FFFF;
defparam prom_inst_27.INIT_RAM_37 = 256'hFFFFE0000007FF71D1FCCFE7F07F1C5FE31FF7DCF9F9CEF83B3FBFFFFFFFFF80;
defparam prom_inst_27.INIT_RAM_38 = 256'h00007FFFBF3F9C6EAE03C383FF79FFFFCFBF9CEF2389C1FFFFFFFFF00007C001;
defparam prom_inst_27.INIT_RAM_39 = 256'hB9EBFEEDC467BC19EFF7BFFFFE7BF8EFF9783F9FFFFFF80000008C000FFFFC00;
defparam prom_inst_27.INIT_RAM_3A = 256'hCC0F3380DE7FBBFF3FE7BF8C6FBB81F9FFFFFFC00000018001FFFFC000001FFF;
defparam prom_inst_27.INIT_RAM_3B = 256'hCE07F0BFF3E6FDE1E0E7B9CFFFFFFFF000000000007FFFFC000001FFF39F3FEE;
defparam prom_inst_27.INIT_RAM_3C = 256'hFF1E0F9E0E06331EFDFFFFFF000000000007FFFF8000001FFF81F3DCE246771B;
defparam prom_inst_27.INIT_RAM_3D = 256'hDFF7EFFFDFBFFFFFFFFFC0003FFFFFFFD0000003FFF83E3E060EF739BEE0FFC1;
defparam prom_inst_27.INIT_RAM_3E = 256'hFFFFFFFFFFFFFE0001FFFFFFF20000007FFFFFF7DFF7CF37DDDEEFFFBFFFFF7F;
defparam prom_inst_27.INIT_RAM_3F = 256'hFFFFFFF0001FFF80000000003FFFFF7FFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_28 (
    .DO({prom_inst_28_dout_w[30:0],prom_inst_28_dout[15]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_32),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_28.READ_MODE = 1'b1;
defparam prom_inst_28.BIT_WIDTH = 1;
defparam prom_inst_28.RESET_MODE = "SYNC";
defparam prom_inst_28.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_04 = 256'hFFFFFFFFFFFC000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_05 = 256'hFFFFE0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_06 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam prom_inst_28.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFF;
defparam prom_inst_28.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0E = 256'hFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0F = 256'hFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_10 = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_28.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFF;
defparam prom_inst_28.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_19 = 256'hFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1A = 256'hF80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001F;
defparam prom_inst_28.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFF;
defparam prom_inst_28.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_23 = 256'hFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_24 = 256'hFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_25 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_28.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFF;
defparam prom_inst_28.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001FFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2D = 256'hFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2E = 256'hFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2F = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_28.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00003FFFF;
defparam prom_inst_28.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_37 = 256'hFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_38 = 256'hFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_28.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FF;
defparam prom_inst_28.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFF;
defparam prom_inst_28.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000003FFFFFFF;
defparam prom_inst_28.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000003FFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFC0000000000000000000000007FFFFFFFFFFFFFFFFFFF;

pROM prom_inst_29 (
    .DO({prom_inst_29_dout_w[30:0],prom_inst_29_dout[15]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_33),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_29.READ_MODE = 1'b1;
defparam prom_inst_29.BIT_WIDTH = 1;
defparam prom_inst_29.RESET_MODE = "SYNC";
defparam prom_inst_29.INIT_RAM_00 = 256'hFFFFFFFFFFFFE0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_01 = 256'hDDEFFFFFFFFFFFFC0001FFF00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_02 = 256'hFFFFFFFFC0001FFFC00000003FFF7FFDC3BF9F97CF93F7BF070C0D93C9B37DB7;
defparam prom_inst_29.INIT_RAM_03 = 256'hFE0001FFFE00000001FFFBDBDFBBF9F7BCFBBF7FFDFEFBDDFBDFBBDBB9DEFFFF;
defparam prom_inst_29.INIT_RAM_04 = 256'hFFF00000000FFFBDBDFDBFAF7BDFFDFFDFDFEFBDDFBDFFBDBB9DEFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_05 = 256'h00007FFBDDDFDDFBFFBD7FDFBDFFFF7BEEFBDFDFDBBBDF7FFFFFFFFFFFE0000F;
defparam prom_inst_29.INIT_RAM_06 = 256'hBDDDFDDFB7FBDFFDFBDFEFF7BEFFDDFDDDDBAFF7FFFFFFFFFFFE0000FFFF8000;
defparam prom_inst_29.INIT_RAM_07 = 256'hFBFDDDBFBFBDFEFF7FEF7ECFDDDDDAEF7FFC0000000FF00007FFF800000003FF;
defparam prom_inst_29.INIT_RAM_08 = 256'hE7FBEFEFF7DEFBE0FDEDDDEEF7FFC00000007F00007FFFC00000001FFBEEFFDD;
defparam prom_inst_29.INIT_RAM_09 = 256'hFFBDFF9EEFFEDDD7EFBFFFFFF00007F00007FFFC00000000FFFEEFFDDFBFC1DD;
defparam prom_inst_29.INIT_RAM_0A = 256'hEEFEF5ED76FBFFFFFF80003F00003FFFE00000000FFDEFDFEDF9BDDDDCFFFEFE;
defparam prom_inst_29.INIT_RAM_0B = 256'hE777BFFFFFFC0003F80003FFFE000000007FDEF7FEFF99DDCDDFFDEFFFFBDF7D;
defparam prom_inst_29.INIT_RAM_0C = 256'hFFFFC0003F80003FFFE000000003FDF7FFEEFBDDEDEDFFDFFF7FBDF7EEEFEF5E;
defparam prom_inst_29.INIT_RAM_0D = 256'h01FC0001FFFF000000003FFF7BFEEEBFDEDEDF7DFFF7FBEF7EEF7EF9EE777BFF;
defparam prom_inst_29.INIT_RAM_0E = 256'h1FFFF000000001FEF79FEEEBEDEDF6E7EEFF7FBEF7F6F7EF9EE773BFFFFFFE00;
defparam prom_inst_29.INIT_RAM_0F = 256'h0000001FFEFDFE75FFDFDF7CFFCFF7FBEFFF6F7E79FEFFB3FFFFFFE0001FC000;
defparam prom_inst_29.INIT_RAM_10 = 256'hFFDFFFFF9FFFFFFF9FF9FFFFFFFFFFFFFFFFFFFE7FFFFFFF0001FC0001FFFF00;
defparam prom_inst_29.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FE0000FFFF000000001;
defparam prom_inst_29.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FE0000FFFF000000000FFFFFFF;
defparam prom_inst_29.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FE00007FFF000000000FFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFC0007F00007FFE0000000007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_15 = 256'hFFFFFFFFFFFFFC0007F00007FFE0000000007FFFFFF5FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_16 = 256'hFFFFFFC0007F00007FFE0000000003FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_17 = 256'h0003F80003FFE0000000003FFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_18 = 256'h003FFC0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_29.INIT_RAM_19 = 256'h000000003E7EF7F0FE7BF7BF03E03F07F83F03E77E0FFDF81FFFFFFFE0003F80;
defparam prom_inst_29.INIT_RAM_1A = 256'h01E7E77E07E73F39F03E03F07F03F03E77E07FCF81FFFFFFFE0001F80003FFC0;
defparam prom_inst_29.INIT_RAM_1B = 256'hE63F73F39FFBFCFE73F39FCFF33FE7FCFF9FFFFFFFE0001FC0001FF800000000;
defparam prom_inst_29.INIT_RAM_1C = 256'h39FFBFCFE79F39FCFF93FF7FCFFDFFFFFFFF0001FC0001FF00000000001F7F37;
defparam prom_inst_29.INIT_RAM_1D = 256'hFE79F39FCFFD3FF7FCFFDFFFFFFFF0000FC0000FE00000000001F7F37EF3F73F;
defparam prom_inst_29.INIT_RAM_1E = 256'hFCFFC3F07FCFC1FFFFFFFF8000FE0000FC00000000001F7F87FFBF61F39FF9FC;
defparam prom_inst_29.INIT_RAM_1F = 256'h07FEFC0FFFFFFFF8000FE00000000000000001F7FC3FF9F61F01FC1FCFE79F99;
defparam prom_inst_29.INIT_RAM_20 = 256'hFFFFFFFF80007E00000000000000000F3F83FF9F29F01F81FCFE7DF81FEFFC3F;
defparam prom_inst_29.INIT_RAM_21 = 256'hFC0007F00000000000000000F3F83FF9F09F9CFF9FCFE7DF81FEFF83FF3FEFFC;
defparam prom_inst_29.INIT_RAM_22 = 256'h00003FFC000000000F3F93FF9F09FBCFFDFEFE7DF9DFEFF9BFF3FEFFCFFFFFFF;
defparam prom_inst_29.INIT_RAM_23 = 256'hF000000000F3F33F79F1DF9CFFDFEFF39F9DFEFF9BFF3FEFFCFFFFFFFFC0003F;
defparam prom_inst_29.INIT_RAM_24 = 256'h000FBF33F31F9DF9CFF9FEFF39F9CFE7F3BFF3FE7FCFFFFFFFFC0003F80003FF;
defparam prom_inst_29.INIT_RAM_25 = 256'hBF03F9CF9CF80FE7F81F9CFE7F39F03E07C0FFFFFFFFE0003F80003FFFC00000;
defparam prom_inst_29.INIT_RAM_26 = 256'hF9EF80FE7FC3F9CFE7E39F03E07C0FFFFFFFFE0001F80003FFFE00000000FBF3;
defparam prom_inst_29.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FC0001FFFF00000000FBE79F83F9C;
defparam prom_inst_29.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0001FC0001FFFF80000000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFF0000FC0000FFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2A = 256'hFFFFFFFFFF8000FE0000FFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2B = 256'hFFF8000FE0000FFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2C = 256'h7E0000FFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2D = 256'hFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_29.INIT_RAM_2E = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007F0000F;
defparam prom_inst_29.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007F0000FFFFF000;
defparam prom_inst_29.INIT_RAM_30 = 256'hE7E07CFC3FEF7F818180FB9CCEF8F07FFFFFFFFC0003F8000FFFFF0000001FFF;
defparam prom_inst_29.INIT_RAM_31 = 256'h99FEF7F81C1C0FB9CE6F8F07FFFFFFFFE0003F8000FFFFF0000001FE773981DF;
defparam prom_inst_29.INIT_RAM_32 = 256'hE7FDF3FB9CF278FF3FFFFFFFFE0001F8000FFFFF0000001FE733981DFE3E07CF;
defparam prom_inst_29.INIT_RAM_33 = 256'hBDCFA787F3FFFFFFFFE0001FC000FFFFF0000003FE73B9F9CFE3EE7C79DFE73F;
defparam prom_inst_29.INIT_RAM_34 = 256'h7F3FFFFFFFFF0001FC000FFFFF0000003FF739BFDCFE1EF7D7FDFE73FF7FCF3F;
defparam prom_inst_29.INIT_RAM_35 = 256'hFFFFF0000FC000FFFFF0000003FF739BF9CFE9E77D3F9FE73FF7FCF3F9DEF879;
defparam prom_inst_29.INIT_RAM_36 = 256'h00FC000FFFFF0000007FF7BDBC1CFEDE0393E1FF73FF7C0FBF9CE7879383FFFF;
defparam prom_inst_29.INIT_RAM_37 = 256'hFFFFE0000007FF3BCBC1EFECF039BC3FF7BFF3E0FBFDCE7879B83FFFFFFFFF00;
defparam prom_inst_29.INIT_RAM_38 = 256'h0000FFF39CBFCEFE4F3399CFFF3BFF3FEF9FDCE79793FBFFFFFFFFF8000FC000;
defparam prom_inst_29.INIT_RAM_39 = 256'h39E3FCE6E0F3381CFFF39FF3FEF9FDCE73381FBFFFFFFFFF800078001FFFFE00;
defparam prom_inst_29.INIT_RAM_3A = 256'h6E077B81CEFF39FFBFEF9FDEE73381FBFFFFFE000000000001FFFFC000000FFF;
defparam prom_inst_29.INIT_RAM_3B = 256'hCCCFF91FFBE079C0E6733BDF9FFFFFE000000000003FFFF8000001FFFB9E3FCE;
defparam prom_inst_29.INIT_RAM_3C = 256'hFFBE07DC0F0F7BBCF9FFFFFFFFFC0003FFFFFFFF0000003FFF99E3E0E4EF73B9;
defparam prom_inst_29.INIT_RAM_3D = 256'hE0F8F7BBEFDFFFFFFFFFE0003FFFFFFFE0000007FFFC1F3C0F0CF33B9CE0FF83;
defparam prom_inst_29.INIT_RAM_3E = 256'hFFFFFFFFFFFFFE0003FFFFFFFC000000FFFFC3FBE0F8FFFBBBEF1FFC7FFBE0FD;
defparam prom_inst_29.INIT_RAM_3F = 256'hFFFFFFE000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_30 (
    .DO({promx9_inst_30_dout_w[26:0],promx9_inst_30_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_35),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_30.READ_MODE = 1'b1;
defparam promx9_inst_30.BIT_WIDTH = 9;
defparam promx9_inst_30.RESET_MODE = "SYNC";
defparam promx9_inst_30.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_05 = 288'h4D9ECF6FCFEC7B3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_06 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_30.INIT_RAM_07 = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D76BB5DAED76BB5DAED76BB5DAED76BB5DA6D369B;
defparam promx9_inst_30.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7D;
defparam promx9_inst_30.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_0E = 288'h4DA6D36DCAE774BADEAF77FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_0F = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6D369B5DAED369B4DA6D369B4DA6D36BB5DAED76BB;
defparam promx9_inst_30.INIT_RAM_10 = 288'hFFFFFFF3E7E26D369B4DA6D369B4DA6D369B4DA6D369B5DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_30.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_17 = 288'hFEFF7FBFDFEFF7FA5D5F4FB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_18 = 288'hFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFD;
defparam promx9_inst_30.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFBFCE26D369B4DA6D369B4DA6D369B4DA6D369BFEFF7FBFDFEFF7FBFD;
defparam promx9_inst_30.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_20 = 288'hFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_21 = 288'hEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDFEFF7FBFDF;
defparam promx9_inst_30.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFF2EA6D369B4DA6D369B4DA6D369B4DA6D369B9F7FFFFFF;
defparam promx9_inst_30.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_2A = 288'hDEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF2ED36BB5DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_30.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_33 = 288'h4DA6D369B7E67FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFD71369B4DA6D369B4DA6D369B;
defparam promx9_inst_30.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_3C = 288'h4DA6D369B4DA6D369B5DAFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA74F69B4DA6D369B;
defparam promx9_inst_30.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_30.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_31 (
    .DO({promx9_inst_31_dout_w[26:0],promx9_inst_31_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_37),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_31.READ_MODE = 1'b1;
defparam promx9_inst_31.BIT_WIDTH = 9;
defparam promx9_inst_31.RESET_MODE = "SYNC";
defparam promx9_inst_31.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_05 = 288'h4DA6D369B4DA6D369B4DA6D369B4DFF7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7DB69B;
defparam promx9_inst_31.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_0E = 288'hFFFFFBA9B4DA6D369B4DA6D369B4DA6D369B4DCF2FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_17 = 288'hFFFFFFFFFFFFFE7C9B4DA6D369B4DA6D369B4DA6D369B5DAEDBDFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFF3F3C4DA6D369B4DA6D369B4DA6D369B4DA6FFBFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBE1D4DA6D369B4DA6D369B4DA6D369B4DA6E399F;
defparam promx9_inst_31.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_31 = 288'h4DA6D36BEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDE6DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_31.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_3A = 288'h4DA6D369B4DA6D373CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9F8E26D369B4DA6D369B;
defparam promx9_inst_31.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_31.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_32 (
    .DO({promx9_inst_32_dout_w[26:0],promx9_inst_32_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_39),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_32.READ_MODE = 1'b1;
defparam promx9_inst_32.BIT_WIDTH = 9;
defparam promx9_inst_32.RESET_MODE = "SYNC";
defparam promx9_inst_32.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_03 = 288'h4DA6D369B4DA6D369B4DA6D369BAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEA6D369B;
defparam promx9_inst_32.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_0C = 288'h8F26D369B4DA6D369B4DA6D369B4DA6D367B1EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_15 = 288'hFFFFFFFFFEFCF1369B4DA6D369B4DA6D369B4DA6D369BAE6FFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFF9F4F69B4DA6D369B4DA6D369B4DA6D369B6DC7BFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7D369B4DA6D369B4DA6D369B4DA6D369B4D977FFFF;
defparam promx9_inst_32.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_2F = 288'h4DDF37FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF389B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_32.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_38 = 288'h4DA6D369B4DB6E7DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3ABB4DA6D369B4DA6D369B;
defparam promx9_inst_32.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_32.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_33 (
    .DO({promx9_inst_33_dout_w[26:0],promx9_inst_33_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_41),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_33.READ_MODE = 1'b1;
defparam promx9_inst_33.BIT_WIDTH = 9;
defparam promx9_inst_33.RESET_MODE = "SYNC";
defparam promx9_inst_33.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_01 = 288'h4DA6D369B4DA6D369B4DA6CBBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBCFC4DA6D369B;
defparam promx9_inst_33.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_0A = 288'h4DA6D369B4DA6D369B4DA6D369B4DA6E39DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFBC;
defparam promx9_inst_33.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_13 = 288'hFFFFFFE7D5DA6D369B4DA6D369B4DA6D369B4DA6CF6FEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFF7E6E26D369B4DA6D369B4DA6D369B4DA6CF7BCFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFCE26D369B4DA6D369B4DA6D369B4DA6D36FCBFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_2D = 288'h4EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6F1ED369B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_33.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_36 = 288'h4DA6D369BCE77FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_33.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_33.INIT_RAM_3F = 288'h4DA6D369B4DA6D369B8DD7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_34 (
    .DO({promx9_inst_34_dout_w[26:0],promx9_inst_34_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_43),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_34.READ_MODE = 1'b1;
defparam promx9_inst_34.BIT_WIDTH = 9;
defparam promx9_inst_34.RESET_MODE = "SYNC";
defparam promx9_inst_34.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF874F69B4DA6D369B;
defparam promx9_inst_34.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_08 = 288'h4DA6D369B4DA6D369B4DA6D369B5DA7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC79769B;
defparam promx9_inst_34.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_11 = 288'hFFEFEF89B4DA6D369B4DA6D369B4DA6D369B4DEF7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_1A = 288'hFFFFFFFFFFFFFCBA9B4DA6D369B4DA6D369B4DA6D369B4DB6F3FFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFDFCDC5DA6D369B4DA6D369B4DA6D369B4DA6CFBFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F5C4DA6D369B4DA6D369B4DA6D369B4DA6E79FF;
defparam promx9_inst_34.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_34 = 288'h4DA6D373EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3D3DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_34.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_3D = 288'h4DA6D369B4DA6D361DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_34.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3E4DA6D369B4DA6D369B;
defparam promx9_inst_34.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_35 (
    .DO({promx9_inst_35_dout_w[26:0],promx9_inst_35_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_45),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_35.READ_MODE = 1'b1;
defparam promx9_inst_35.BIT_WIDTH = 9;
defparam promx9_inst_35.RESET_MODE = "SYNC";
defparam promx9_inst_35.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_06 = 288'h4DA6D369B4DA6D369B5DA6D371CDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8E26D369B;
defparam promx9_inst_35.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_0F = 288'h7F26D369B4DA6D369B4DA6D369B4DA6D36DB7F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_18 = 288'hFFFFFFFFFDFCF1369B4DA6D369B4DA6D369B4DA6D369B0EFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFF975369B4DA6D369B4DA6D369B4DA6D369BAE67FFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD79F89B4DA6D369B4DA6D369B4DA6D369B5DC7BFFFF;
defparam promx9_inst_35.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_32 = 288'h3D877FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FBA9B4DA6D369B4DA6D369B4DA6D369B;
defparam promx9_inst_35.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_3B = 288'h4DA6D369B4DBEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFCBB5DA6D369B4DA6D369B;
defparam promx9_inst_35.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_35.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_36 (
    .DO({promx9_inst_36_dout_w[26:0],promx9_inst_36_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_47),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_36.READ_MODE = 1'b1;
defparam promx9_inst_36.BIT_WIDTH = 9;
defparam promx9_inst_36.RESET_MODE = "SYNC";
defparam promx9_inst_36.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_02 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_04 = 288'h4DA6D369B4DA6D369B4DA6DBDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F9C4DA6D369B;
defparam promx9_inst_36.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_0B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_0D = 288'h5DA6D369B4DA6D369B4DA6D369B4DA6EF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDE;
defparam promx9_inst_36.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_14 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_16 = 288'hFFFFFFFFFBE26D369B4DA6D369B4DA6D369B4DA6CF79FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFAFAED369B4DA6D369B4DA6D369B4DA6D367DFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFEF875769B4DA6D369B4DA6D369B4DA6D379CDFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_30 = 288'h9F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFA789B4DA6D369B4DA6D369B4DA6D36FC;
defparam promx9_inst_36.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_37 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_39 = 288'h4DA6D36BB4F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7CBABB4DA6D369B4DA6D369B;
defparam promx9_inst_36.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_36.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROMX9 promx9_inst_37 (
    .DO({promx9_inst_37_dout_w[26:0],promx9_inst_37_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_49),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam promx9_inst_37.READ_MODE = 1'b1;
defparam promx9_inst_37.BIT_WIDTH = 9;
defparam promx9_inst_37.RESET_MODE = "SYNC";
defparam promx9_inst_37.INIT_RAM_00 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_01 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_02 = 288'h4DA6D369B4DA6D369BCEF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_03 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF3C3DAED369B;
defparam promx9_inst_37.INIT_RAM_04 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_05 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_06 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_07 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_08 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_09 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_0A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_0B = 288'h8D9ED369B4DA6D369B4DA6D369B5DE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_0C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F;
defparam promx9_inst_37.INIT_RAM_0D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_0E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_0F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_10 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_11 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_12 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_13 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_14 = 288'hFFFFFFFFF4EBF1369B4DA6D369B4DA6D369B4D977FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_15 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_16 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_17 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_18 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_19 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_1A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_1B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_1C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_1D = 288'hFFFFFFFFFFFFFFFFFFDF8F5F87B4DA6D369B4DA6D369B4DCF3BFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_1E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_1F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_20 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_21 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_22 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_23 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_24 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_25 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_26 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFBABB4DA6D369B4DA6D369B4D9EE7DFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_27 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_28 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_29 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_2A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_2B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_2C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_2D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_2E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_2F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3DA6D369B4DA6D369B4DA6FBBFF;
defparam promx9_inst_37.INIT_RAM_30 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_31 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_32 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_33 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_34 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_35 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_36 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_37 = 288'h4DA6E397FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_38 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7E4F3F0F69B4DA6D369B;
defparam promx9_inst_37.INIT_RAM_39 = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_3A = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_3B = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_3C = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_3D = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_3E = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam promx9_inst_37.INIT_RAM_3F = 288'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_38 (
    .DO({prom_inst_38_dout_w[30:0],prom_inst_38_dout[9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_38.READ_MODE = 1'b1;
defparam prom_inst_38.BIT_WIDTH = 1;
defparam prom_inst_38.RESET_MODE = "SYNC";
defparam prom_inst_38.INIT_RAM_00 = 256'h000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_01 = 256'h0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_02 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam prom_inst_38.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000;
defparam prom_inst_38.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_09 = 256'hFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0A = 256'hFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001F;
defparam prom_inst_38.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFF;
defparam prom_inst_38.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_13 = 256'hFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_14 = 256'hFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_15 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_38.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFF;
defparam prom_inst_38.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_1D = 256'hFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_1E = 256'hFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_1F = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_38.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFF;
defparam prom_inst_38.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_27 = 256'hFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_28 = 256'hFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_29 = 256'h8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFF;
defparam prom_inst_38.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_32 = 256'hFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_33 = 256'hFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000F;
defparam prom_inst_38.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFF;
defparam prom_inst_38.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3C = 256'hFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3D = 256'hFFFFE001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3E = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;

pROM prom_inst_39 (
    .DO({prom_inst_39_dout_w[30:0],prom_inst_39_dout[10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_39.READ_MODE = 1'b1;
defparam prom_inst_39.BIT_WIDTH = 1;
defparam prom_inst_39.RESET_MODE = "SYNC";
defparam prom_inst_39.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_40 (
    .DO({prom_inst_40_dout_w[30:0],prom_inst_40_dout[11]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_40.READ_MODE = 1'b1;
defparam prom_inst_40.BIT_WIDTH = 1;
defparam prom_inst_40.RESET_MODE = "SYNC";
defparam prom_inst_40.INIT_RAM_00 = 256'h0000000C0000000005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_01 = 256'h00000000153FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_40.INIT_RAM_02 = 256'h00DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000800;
defparam prom_inst_40.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80008000000000;
defparam prom_inst_40.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000707FFC000F9FFFFFF;
defparam prom_inst_40.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFC0005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_09 = 256'hFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0A = 256'hFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0003F;
defparam prom_inst_40.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0002FFFFFFFF;
defparam prom_inst_40.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00017FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_13 = 256'hFFFFFFFFFF8000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_14 = 256'hFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_15 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_40.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFF;
defparam prom_inst_40.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0003FFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1D = 256'hFFFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1E = 256'hFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1F = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_40.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA000FFFFF;
defparam prom_inst_40.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0005FFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0005FFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_27 = 256'hFFFFFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_28 = 256'hFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_29 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFF;
defparam prom_inst_40.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_32 = 256'hFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_33 = 256'hFF4000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4000F;
defparam prom_inst_40.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA000FFFFFFFF;
defparam prom_inst_40.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9001FFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD000BFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF4003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFA005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3C = 256'hFFFFFFFFFFFE003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3D = 256'hFFFFE001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3E = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;

pROM prom_inst_41 (
    .DO({prom_inst_41_dout_w[30:0],prom_inst_41_dout[12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_41.READ_MODE = 1'b1;
defparam prom_inst_41.BIT_WIDTH = 1;
defparam prom_inst_41.RESET_MODE = "SYNC";
defparam prom_inst_41.INIT_RAM_00 = 256'h0001FFF0000000000DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_01 = 256'h0000000010FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_02 = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000;
defparam prom_inst_41.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000;
defparam prom_inst_41.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007F8003FFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_09 = 256'hFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0A = 256'hFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0001F;
defparam prom_inst_41.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFF;
defparam prom_inst_41.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8000FFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFF4000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_13 = 256'hFFFFFFFFFFC000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_14 = 256'hFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_15 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_41.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0005FFFFFF;
defparam prom_inst_41.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1D = 256'hFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1E = 256'hFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1F = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_41.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0007FFFF;
defparam prom_inst_41.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0005FFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFD0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_27 = 256'hFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_28 = 256'hFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_29 = 256'h8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4000FFF;
defparam prom_inst_41.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFD0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_32 = 256'hFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_33 = 256'hFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80017;
defparam prom_inst_41.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFF;
defparam prom_inst_41.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF2007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3C = 256'hFFFFFFFFFFFB001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3D = 256'hFFFFF003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3E = 256'h2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;

pROM prom_inst_42 (
    .DO({prom_inst_42_dout_w[30:0],prom_inst_42_dout[13]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_42.READ_MODE = 1'b1;
defparam prom_inst_42.BIT_WIDTH = 1;
defparam prom_inst_42.RESET_MODE = "SYNC";
defparam prom_inst_42.INIT_RAM_00 = 256'h00000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_01 = 256'h00000000057FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_42.INIT_RAM_02 = 256'hFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8000000;
defparam prom_inst_42.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_09 = 256'hFFFFFFFFE0005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0A = 256'hFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0003F;
defparam prom_inst_42.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFF;
defparam prom_inst_42.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_13 = 256'hFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_14 = 256'hFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_15 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_42.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFF;
defparam prom_inst_42.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0001FFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1D = 256'hFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1E = 256'hFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1F = 256'h00BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_42.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFF;
defparam prom_inst_42.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_27 = 256'hFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_28 = 256'hFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_29 = 256'h8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFF;
defparam prom_inst_42.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0007FFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_32 = 256'hFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_33 = 256'hFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000F;
defparam prom_inst_42.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0017FFFFFFF;
defparam prom_inst_42.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8003FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3C = 256'hFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3D = 256'hFFFFF003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3E = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE40;

pROM prom_inst_43 (
    .DO({prom_inst_43_dout_w[30:0],prom_inst_43_dout[14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_43.READ_MODE = 1'b1;
defparam prom_inst_43.BIT_WIDTH = 1;
defparam prom_inst_43.RESET_MODE = "SYNC";
defparam prom_inst_43.INIT_RAM_00 = 256'h00000000000000000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_01 = 256'h000000000CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_43.INIT_RAM_02 = 256'hFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam prom_inst_43.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_09 = 256'hFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0A = 256'hFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003F;
defparam prom_inst_43.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFF;
defparam prom_inst_43.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_13 = 256'hFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_14 = 256'hFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_15 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_43.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFF;
defparam prom_inst_43.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1D = 256'hFFFFFFFFFFFF00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1E = 256'hFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1F = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_43.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFF;
defparam prom_inst_43.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_27 = 256'hFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_28 = 256'hFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_29 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFF;
defparam prom_inst_43.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_32 = 256'hFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_33 = 256'hFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001F;
defparam prom_inst_43.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFF;
defparam prom_inst_43.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3C = 256'hFFFFFFFFFFFE003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3D = 256'hFFFFF003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3E = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;

pROM prom_inst_44 (
    .DO({prom_inst_44_dout_w[30:0],prom_inst_44_dout[15]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_50),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_44.READ_MODE = 1'b1;
defparam prom_inst_44.BIT_WIDTH = 1;
defparam prom_inst_44.RESET_MODE = "SYNC";
defparam prom_inst_44.INIT_RAM_00 = 256'h000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_01 = 256'h0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_02 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam prom_inst_44.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000;
defparam prom_inst_44.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_09 = 256'hFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0A = 256'hFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001F;
defparam prom_inst_44.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFF;
defparam prom_inst_44.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_13 = 256'hFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_14 = 256'hFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_15 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam prom_inst_44.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFF;
defparam prom_inst_44.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1D = 256'hFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1E = 256'hFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1F = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam prom_inst_44.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFF;
defparam prom_inst_44.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_27 = 256'hFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_28 = 256'hFFFFFFF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_29 = 256'h8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FF;
defparam prom_inst_44.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_32 = 256'hFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_33 = 256'hFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000F;
defparam prom_inst_44.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFF;
defparam prom_inst_44.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3C = 256'hFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3D = 256'hFFFFE001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3E = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;

pROM prom_inst_45 (
    .DO({prom_inst_45_dout_w[15:0],prom_inst_45_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_52),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_45.READ_MODE = 1'b1;
defparam prom_inst_45.BIT_WIDTH = 16;
defparam prom_inst_45.RESET_MODE = "SYNC";
defparam prom_inst_45.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_01 = 256'h049B047B049B049B049B049B0CBBA6BEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE79F9EBE65DC24FC;
defparam prom_inst_45.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_13 = 256'hFFFFFFFFCF5E863D4D9C3D3C351C24FC1CDB24FC2D1C8E7DFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_24 = 256'hF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFBFBEDE9E7E75DD557C6DBD8E3EBEFE;
defparam prom_inst_45.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_5 (
  .Q(dff_q_5),
  .D(dff_q_4),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_6 (
  .Q(dff_q_6),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_7 (
  .Q(dff_q_7),
  .D(dff_q_6),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_8 (
  .Q(dff_q_8),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_9 (
  .Q(dff_q_9),
  .D(dff_q_8),
  .CLK(clk),
  .CE(oce)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(promx9_inst_0_dout[0]),
  .I1(promx9_inst_1_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(promx9_inst_2_dout[0]),
  .I1(promx9_inst_3_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(promx9_inst_4_dout[0]),
  .I1(promx9_inst_5_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(promx9_inst_6_dout[0]),
  .I1(promx9_inst_7_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(promx9_inst_8_dout[0]),
  .I1(promx9_inst_9_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(promx9_inst_10_dout[0]),
  .I1(promx9_inst_11_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(promx9_inst_12_dout[0]),
  .I1(promx9_inst_13_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(promx9_inst_14_dout[0]),
  .I1(promx9_inst_15_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(promx9_inst_30_dout[0]),
  .I1(promx9_inst_31_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(promx9_inst_32_dout[0]),
  .I1(promx9_inst_33_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(promx9_inst_34_dout[0]),
  .I1(promx9_inst_35_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(promx9_inst_36_dout[0]),
  .I1(promx9_inst_37_dout[0]),
  .S0(dff_q_9)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(dff_q_7)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_27),
  .I1(mux_o_28),
  .S0(dff_q_7)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_29),
  .I1(mux_o_30),
  .S0(dff_q_7)
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_31),
  .I1(mux_o_32),
  .S0(dff_q_7)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(dff_q_7)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_7)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(dff_q_5)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(dff_q_5)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_5)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_3)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_47),
  .I1(prom_inst_45_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_51 (
  .O(dout[0]),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_1)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(promx9_inst_0_dout[1]),
  .I1(promx9_inst_1_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(promx9_inst_2_dout[1]),
  .I1(promx9_inst_3_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(promx9_inst_4_dout[1]),
  .I1(promx9_inst_5_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(promx9_inst_6_dout[1]),
  .I1(promx9_inst_7_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(promx9_inst_8_dout[1]),
  .I1(promx9_inst_9_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(promx9_inst_10_dout[1]),
  .I1(promx9_inst_11_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(promx9_inst_12_dout[1]),
  .I1(promx9_inst_13_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(promx9_inst_14_dout[1]),
  .I1(promx9_inst_15_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(promx9_inst_30_dout[1]),
  .I1(promx9_inst_31_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(promx9_inst_32_dout[1]),
  .I1(promx9_inst_33_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(promx9_inst_34_dout[1]),
  .I1(promx9_inst_35_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(promx9_inst_36_dout[1]),
  .I1(promx9_inst_37_dout[1]),
  .S0(dff_q_9)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_7)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_7)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_7)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(dff_q_7)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_7)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(dff_q_7)
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(dff_q_5)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(dff_q_5)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(dff_q_5)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_97),
  .I1(mux_o_98),
  .S0(dff_q_3)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_99),
  .I1(prom_inst_45_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_103 (
  .O(dout[1]),
  .I0(mux_o_101),
  .I1(mux_o_102),
  .S0(dff_q_1)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(promx9_inst_0_dout[2]),
  .I1(promx9_inst_1_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(promx9_inst_2_dout[2]),
  .I1(promx9_inst_3_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(promx9_inst_4_dout[2]),
  .I1(promx9_inst_5_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(promx9_inst_6_dout[2]),
  .I1(promx9_inst_7_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(promx9_inst_8_dout[2]),
  .I1(promx9_inst_9_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(promx9_inst_10_dout[2]),
  .I1(promx9_inst_11_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(promx9_inst_12_dout[2]),
  .I1(promx9_inst_13_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(promx9_inst_14_dout[2]),
  .I1(promx9_inst_15_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(promx9_inst_30_dout[2]),
  .I1(promx9_inst_31_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(promx9_inst_32_dout[2]),
  .I1(promx9_inst_33_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(promx9_inst_34_dout[2]),
  .I1(promx9_inst_35_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(promx9_inst_36_dout[2]),
  .I1(promx9_inst_37_dout[2]),
  .S0(dff_q_9)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(mux_o_129),
  .I1(mux_o_130),
  .S0(dff_q_7)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_131),
  .I1(mux_o_132),
  .S0(dff_q_7)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(dff_q_7)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_7)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_7)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(dff_q_7)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(dff_q_5)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(dff_q_5)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(dff_q_5)
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(mux_o_149),
  .I1(mux_o_150),
  .S0(dff_q_3)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(mux_o_151),
  .I1(prom_inst_45_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_155 (
  .O(dout[2]),
  .I0(mux_o_153),
  .I1(mux_o_154),
  .S0(dff_q_1)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(promx9_inst_0_dout[3]),
  .I1(promx9_inst_1_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(promx9_inst_2_dout[3]),
  .I1(promx9_inst_3_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(promx9_inst_4_dout[3]),
  .I1(promx9_inst_5_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(promx9_inst_6_dout[3]),
  .I1(promx9_inst_7_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(promx9_inst_8_dout[3]),
  .I1(promx9_inst_9_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(promx9_inst_10_dout[3]),
  .I1(promx9_inst_11_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(promx9_inst_12_dout[3]),
  .I1(promx9_inst_13_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(promx9_inst_14_dout[3]),
  .I1(promx9_inst_15_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(promx9_inst_30_dout[3]),
  .I1(promx9_inst_31_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(promx9_inst_32_dout[3]),
  .I1(promx9_inst_33_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(promx9_inst_34_dout[3]),
  .I1(promx9_inst_35_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(promx9_inst_36_dout[3]),
  .I1(promx9_inst_37_dout[3]),
  .S0(dff_q_9)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_7)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(dff_q_7)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(mux_o_185),
  .I1(mux_o_186),
  .S0(dff_q_7)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(mux_o_187),
  .I1(mux_o_188),
  .S0(dff_q_7)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(dff_q_7)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(dff_q_7)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(dff_q_5)
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_5)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_5)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(dff_q_3)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_203),
  .I1(prom_inst_45_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_207 (
  .O(dout[3]),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_1)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(promx9_inst_0_dout[4]),
  .I1(promx9_inst_1_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(promx9_inst_2_dout[4]),
  .I1(promx9_inst_3_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(promx9_inst_4_dout[4]),
  .I1(promx9_inst_5_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(promx9_inst_6_dout[4]),
  .I1(promx9_inst_7_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(promx9_inst_8_dout[4]),
  .I1(promx9_inst_9_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(promx9_inst_10_dout[4]),
  .I1(promx9_inst_11_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(promx9_inst_12_dout[4]),
  .I1(promx9_inst_13_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(promx9_inst_14_dout[4]),
  .I1(promx9_inst_15_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(promx9_inst_30_dout[4]),
  .I1(promx9_inst_31_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(promx9_inst_32_dout[4]),
  .I1(promx9_inst_33_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(promx9_inst_34_dout[4]),
  .I1(promx9_inst_35_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(promx9_inst_36_dout[4]),
  .I1(promx9_inst_37_dout[4]),
  .S0(dff_q_9)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_7)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_7)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(dff_q_7)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(dff_q_7)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(dff_q_7)
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(dff_q_7)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(mux_o_246),
  .I1(mux_o_247),
  .S0(dff_q_5)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(dff_q_5)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(dff_q_5)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(mux_o_253),
  .I1(mux_o_254),
  .S0(dff_q_3)
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(mux_o_255),
  .I1(prom_inst_45_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_259 (
  .O(dout[4]),
  .I0(mux_o_257),
  .I1(mux_o_258),
  .S0(dff_q_1)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(promx9_inst_0_dout[5]),
  .I1(promx9_inst_1_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(promx9_inst_2_dout[5]),
  .I1(promx9_inst_3_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(promx9_inst_4_dout[5]),
  .I1(promx9_inst_5_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(promx9_inst_6_dout[5]),
  .I1(promx9_inst_7_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(promx9_inst_8_dout[5]),
  .I1(promx9_inst_9_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(promx9_inst_10_dout[5]),
  .I1(promx9_inst_11_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(promx9_inst_12_dout[5]),
  .I1(promx9_inst_13_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(promx9_inst_14_dout[5]),
  .I1(promx9_inst_15_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(promx9_inst_30_dout[5]),
  .I1(promx9_inst_31_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(promx9_inst_32_dout[5]),
  .I1(promx9_inst_33_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(promx9_inst_34_dout[5]),
  .I1(promx9_inst_35_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(promx9_inst_36_dout[5]),
  .I1(promx9_inst_37_dout[5]),
  .S0(dff_q_9)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_285),
  .I1(mux_o_286),
  .S0(dff_q_7)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_7)
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_7)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_7)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(mux_o_293),
  .I1(mux_o_294),
  .S0(dff_q_7)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_295),
  .I1(mux_o_296),
  .S0(dff_q_7)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(dff_q_5)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(dff_q_5)
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(dff_q_5)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(dff_q_3)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(mux_o_307),
  .I1(prom_inst_45_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_311 (
  .O(dout[5]),
  .I0(mux_o_309),
  .I1(mux_o_310),
  .S0(dff_q_1)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(promx9_inst_0_dout[6]),
  .I1(promx9_inst_1_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(promx9_inst_2_dout[6]),
  .I1(promx9_inst_3_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(promx9_inst_4_dout[6]),
  .I1(promx9_inst_5_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(promx9_inst_6_dout[6]),
  .I1(promx9_inst_7_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(promx9_inst_8_dout[6]),
  .I1(promx9_inst_9_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(promx9_inst_10_dout[6]),
  .I1(promx9_inst_11_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(promx9_inst_12_dout[6]),
  .I1(promx9_inst_13_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(promx9_inst_14_dout[6]),
  .I1(promx9_inst_15_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(promx9_inst_30_dout[6]),
  .I1(promx9_inst_31_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(promx9_inst_32_dout[6]),
  .I1(promx9_inst_33_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(promx9_inst_34_dout[6]),
  .I1(promx9_inst_35_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(promx9_inst_36_dout[6]),
  .I1(promx9_inst_37_dout[6]),
  .S0(dff_q_9)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(mux_o_337),
  .I1(mux_o_338),
  .S0(dff_q_7)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(mux_o_339),
  .I1(mux_o_340),
  .S0(dff_q_7)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(mux_o_341),
  .I1(mux_o_342),
  .S0(dff_q_7)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(dff_q_7)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_7)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_7)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(dff_q_5)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(dff_q_5)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(dff_q_5)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_3)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_359),
  .I1(prom_inst_45_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_363 (
  .O(dout[6]),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(dff_q_1)
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(promx9_inst_0_dout[7]),
  .I1(promx9_inst_1_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(promx9_inst_2_dout[7]),
  .I1(promx9_inst_3_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(promx9_inst_4_dout[7]),
  .I1(promx9_inst_5_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(promx9_inst_6_dout[7]),
  .I1(promx9_inst_7_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(promx9_inst_8_dout[7]),
  .I1(promx9_inst_9_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(promx9_inst_10_dout[7]),
  .I1(promx9_inst_11_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(promx9_inst_12_dout[7]),
  .I1(promx9_inst_13_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(promx9_inst_14_dout[7]),
  .I1(promx9_inst_15_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(promx9_inst_30_dout[7]),
  .I1(promx9_inst_31_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(promx9_inst_32_dout[7]),
  .I1(promx9_inst_33_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(promx9_inst_34_dout[7]),
  .I1(promx9_inst_35_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(promx9_inst_36_dout[7]),
  .I1(promx9_inst_37_dout[7]),
  .S0(dff_q_9)
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(mux_o_389),
  .I1(mux_o_390),
  .S0(dff_q_7)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(mux_o_391),
  .I1(mux_o_392),
  .S0(dff_q_7)
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(mux_o_393),
  .I1(mux_o_394),
  .S0(dff_q_7)
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(mux_o_395),
  .I1(mux_o_396),
  .S0(dff_q_7)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(mux_o_397),
  .I1(mux_o_398),
  .S0(dff_q_7)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(mux_o_399),
  .I1(mux_o_400),
  .S0(dff_q_7)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(dff_q_5)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(mux_o_404),
  .I1(mux_o_405),
  .S0(dff_q_5)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(mux_o_406),
  .I1(mux_o_407),
  .S0(dff_q_5)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(dff_q_3)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_411),
  .I1(prom_inst_45_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_415 (
  .O(dout[7]),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_1)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(promx9_inst_0_dout[8]),
  .I1(promx9_inst_1_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(promx9_inst_2_dout[8]),
  .I1(promx9_inst_3_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(promx9_inst_4_dout[8]),
  .I1(promx9_inst_5_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(promx9_inst_6_dout[8]),
  .I1(promx9_inst_7_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(promx9_inst_8_dout[8]),
  .I1(promx9_inst_9_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(promx9_inst_10_dout[8]),
  .I1(promx9_inst_11_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_447 (
  .O(mux_o_447),
  .I0(promx9_inst_12_dout[8]),
  .I1(promx9_inst_13_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_448 (
  .O(mux_o_448),
  .I0(promx9_inst_14_dout[8]),
  .I1(promx9_inst_15_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_449 (
  .O(mux_o_449),
  .I0(promx9_inst_30_dout[8]),
  .I1(promx9_inst_31_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_450 (
  .O(mux_o_450),
  .I0(promx9_inst_32_dout[8]),
  .I1(promx9_inst_33_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_451 (
  .O(mux_o_451),
  .I0(promx9_inst_34_dout[8]),
  .I1(promx9_inst_35_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_452 (
  .O(mux_o_452),
  .I0(promx9_inst_36_dout[8]),
  .I1(promx9_inst_37_dout[8]),
  .S0(dff_q_9)
);
MUX2 mux_inst_454 (
  .O(mux_o_454),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(dff_q_7)
);
MUX2 mux_inst_455 (
  .O(mux_o_455),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(dff_q_7)
);
MUX2 mux_inst_456 (
  .O(mux_o_456),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(dff_q_7)
);
MUX2 mux_inst_457 (
  .O(mux_o_457),
  .I0(mux_o_447),
  .I1(mux_o_448),
  .S0(dff_q_7)
);
MUX2 mux_inst_458 (
  .O(mux_o_458),
  .I0(mux_o_449),
  .I1(mux_o_450),
  .S0(dff_q_7)
);
MUX2 mux_inst_459 (
  .O(mux_o_459),
  .I0(mux_o_451),
  .I1(mux_o_452),
  .S0(dff_q_7)
);
MUX2 mux_inst_461 (
  .O(mux_o_461),
  .I0(mux_o_454),
  .I1(mux_o_455),
  .S0(dff_q_5)
);
MUX2 mux_inst_462 (
  .O(mux_o_462),
  .I0(mux_o_456),
  .I1(mux_o_457),
  .S0(dff_q_5)
);
MUX2 mux_inst_463 (
  .O(mux_o_463),
  .I0(mux_o_458),
  .I1(mux_o_459),
  .S0(dff_q_5)
);
MUX2 mux_inst_465 (
  .O(mux_o_465),
  .I0(mux_o_461),
  .I1(mux_o_462),
  .S0(dff_q_3)
);
MUX2 mux_inst_466 (
  .O(mux_o_466),
  .I0(mux_o_463),
  .I1(prom_inst_45_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_467 (
  .O(dout[8]),
  .I0(mux_o_465),
  .I1(mux_o_466),
  .S0(dff_q_1)
);
MUX2 mux_inst_484 (
  .O(mux_o_484),
  .I0(prom_inst_16_dout[9]),
  .I1(prom_inst_17_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_485 (
  .O(mux_o_485),
  .I0(prom_inst_38_dout[9]),
  .I1(prom_inst_45_dout[9]),
  .S0(dff_q_3)
);
MUX2 mux_inst_486 (
  .O(dout[9]),
  .I0(mux_o_484),
  .I1(mux_o_485),
  .S0(dff_q_1)
);
MUX2 mux_inst_503 (
  .O(mux_o_503),
  .I0(prom_inst_18_dout[10]),
  .I1(prom_inst_19_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_504 (
  .O(mux_o_504),
  .I0(prom_inst_39_dout[10]),
  .I1(prom_inst_45_dout[10]),
  .S0(dff_q_3)
);
MUX2 mux_inst_505 (
  .O(dout[10]),
  .I0(mux_o_503),
  .I1(mux_o_504),
  .S0(dff_q_1)
);
MUX2 mux_inst_522 (
  .O(mux_o_522),
  .I0(prom_inst_20_dout[11]),
  .I1(prom_inst_21_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_523 (
  .O(mux_o_523),
  .I0(prom_inst_40_dout[11]),
  .I1(prom_inst_45_dout[11]),
  .S0(dff_q_3)
);
MUX2 mux_inst_524 (
  .O(dout[11]),
  .I0(mux_o_522),
  .I1(mux_o_523),
  .S0(dff_q_1)
);
MUX2 mux_inst_541 (
  .O(mux_o_541),
  .I0(prom_inst_22_dout[12]),
  .I1(prom_inst_23_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_542 (
  .O(mux_o_542),
  .I0(prom_inst_41_dout[12]),
  .I1(prom_inst_45_dout[12]),
  .S0(dff_q_3)
);
MUX2 mux_inst_543 (
  .O(dout[12]),
  .I0(mux_o_541),
  .I1(mux_o_542),
  .S0(dff_q_1)
);
MUX2 mux_inst_560 (
  .O(mux_o_560),
  .I0(prom_inst_24_dout[13]),
  .I1(prom_inst_25_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_561 (
  .O(mux_o_561),
  .I0(prom_inst_42_dout[13]),
  .I1(prom_inst_45_dout[13]),
  .S0(dff_q_3)
);
MUX2 mux_inst_562 (
  .O(dout[13]),
  .I0(mux_o_560),
  .I1(mux_o_561),
  .S0(dff_q_1)
);
MUX2 mux_inst_579 (
  .O(mux_o_579),
  .I0(prom_inst_26_dout[14]),
  .I1(prom_inst_27_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_580 (
  .O(mux_o_580),
  .I0(prom_inst_43_dout[14]),
  .I1(prom_inst_45_dout[14]),
  .S0(dff_q_3)
);
MUX2 mux_inst_581 (
  .O(dout[14]),
  .I0(mux_o_579),
  .I1(mux_o_580),
  .S0(dff_q_1)
);
MUX2 mux_inst_598 (
  .O(mux_o_598),
  .I0(prom_inst_28_dout[15]),
  .I1(prom_inst_29_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_599 (
  .O(mux_o_599),
  .I0(prom_inst_44_dout[15]),
  .I1(prom_inst_45_dout[15]),
  .S0(dff_q_3)
);
MUX2 mux_inst_600 (
  .O(dout[15]),
  .I0(mux_o_598),
  .I1(mux_o_599),
  .S0(dff_q_1)
);
endmodule //Gowin_pROM2
