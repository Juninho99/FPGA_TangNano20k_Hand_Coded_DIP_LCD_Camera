//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Tue Aug 08 19:44:44 2023

module Gowin_SDPB3 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb); //630x390+1

output [0:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [17:0] ada;
input [0:0] din;
input [17:0] adb;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [0:0] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [0:0] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [0:0] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [0:0] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [0:0] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [0:0] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [0:0] sdpb_inst_7_dout;
wire [30:0] sdpb_inst_8_dout_w;
wire [0:0] sdpb_inst_8_dout;
wire [30:0] sdpb_inst_9_dout_w;
wire [0:0] sdpb_inst_9_dout;
wire [30:0] sdpb_inst_10_dout_w;
wire [0:0] sdpb_inst_10_dout;
wire [30:0] sdpb_inst_11_dout_w;
wire [0:0] sdpb_inst_11_dout;
wire [30:0] sdpb_inst_12_dout_w;
wire [0:0] sdpb_inst_12_dout;
wire [30:0] sdpb_inst_13_dout_w;
wire [0:0] sdpb_inst_13_dout;
wire [30:0] sdpb_inst_14_dout_w;
wire [0:0] sdpb_inst_14_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_8.INIT = 16'h0100;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_9.INIT = 16'h0200;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_10.INIT = 16'h0400;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_11.INIT = 16'h0800;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_12.INIT = 16'h1000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_13.INIT = 16'h2000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_14.INIT = 16'h4000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_15.INIT = 16'h0001;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_16.INIT = 16'h0002;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_17.INIT = 16'h0004;
LUT4 lut_inst_18 (
  .F(lut_f_18),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_18.INIT = 16'h0008;
LUT4 lut_inst_19 (
  .F(lut_f_19),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_19.INIT = 16'h0010;
LUT4 lut_inst_20 (
  .F(lut_f_20),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_20.INIT = 16'h0020;
LUT4 lut_inst_21 (
  .F(lut_f_21),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_21.INIT = 16'h0040;
LUT4 lut_inst_22 (
  .F(lut_f_22),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_22.INIT = 16'h0080;
LUT4 lut_inst_23 (
  .F(lut_f_23),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_23.INIT = 16'h0100;
LUT4 lut_inst_24 (
  .F(lut_f_24),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_24.INIT = 16'h0200;
LUT4 lut_inst_25 (
  .F(lut_f_25),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_25.INIT = 16'h0400;
LUT4 lut_inst_26 (
  .F(lut_f_26),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_26.INIT = 16'h0800;
LUT4 lut_inst_27 (
  .F(lut_f_27),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_27.INIT = 16'h1000;
LUT4 lut_inst_28 (
  .F(lut_f_28),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_28.INIT = 16'h2000;
LUT4 lut_inst_29 (
  .F(lut_f_29),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_29.INIT = 16'h4000;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_15}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00007FFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000003FFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFF;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000007FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hFFFFF80000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000001FFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000007FFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFC00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000003FFFFF;
defparam sdpb_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFE000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000001;
defparam sdpb_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam sdpb_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_36 = 256'hFC000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000007FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3B = 256'hFFFFFFE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_16}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFF000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000001FFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFF8000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000FFF;
defparam sdpb_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFF8000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam sdpb_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam sdpb_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_16 = 256'hFFF8000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1B = 256'hFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFF;
defparam sdpb_inst_1.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFE0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000F;
defparam sdpb_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam sdpb_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_36 = 256'hFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_17}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003FFFF;
defparam sdpb_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000;
defparam sdpb_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam sdpb_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_11 = 256'hFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_16 = 256'hFFFFFFC0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1B = 256'hFFFFFFFFFFFE0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000FFF;
defparam sdpb_inst_2.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_27 = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000;
defparam sdpb_inst_2.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2C = 256'h00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam sdpb_inst_2.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_31 = 256'hFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_36 = 256'hFFFFFFFF8000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003FFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFF;
defparam sdpb_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_18}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001F;
defparam sdpb_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000;
defparam sdpb_inst_3.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0C = 256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_3.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_11 = 256'hFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_16 = 256'hFFFFFFFFFE0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFF;
defparam sdpb_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000;
defparam sdpb_inst_3.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_27 = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam sdpb_inst_3.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2C = 256'hF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_31 = 256'hFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_36 = 256'hFFFFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000001FFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFF;
defparam sdpb_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_19}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFE0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_02 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000;
defparam sdpb_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_07 = 256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000001FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0C = 256'hFFE0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_11 = 256'hFFFFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000007FFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_16 = 256'hFFFFFFFFFFFFF8000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFF;
defparam sdpb_inst_4.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFF8000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003F;
defparam sdpb_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_22 = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000;
defparam sdpb_inst_4.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_27 = 256'h000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam sdpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2A = 256'hFFFFFFFFFFFFE00000000000000000000000000000000000000000000000001F;
defparam sdpb_inst_4.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2C = 256'h00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000;
defparam sdpb_inst_4.INIT_RAM_2E = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_31 = 256'h000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000;
defparam sdpb_inst_4.INIT_RAM_33 = 256'h0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_36 = 256'h000000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000;
defparam sdpb_inst_4.INIT_RAM_38 = 256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3B = 256'h000000000000000000000000000000000000000000000000000001FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sdpb_inst_4.INIT_RAM_3D = 256'h0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3E = 256'hFFFFFFFFFF7FFFFFFFEFFEFFFFFFFFFFF8000000000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFDFFFFFFDFFFFFDFFF7FFE3FFFFDFFDFFFFBFFFFBFF9FFDFB;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_20}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b0;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'hFFFF00000000000000000000000000000000000000000000000000000001FFFF;
defparam sdpb_inst_5.INIT_RAM_01 = 256'h3FF0FFF007FFF3FF3FF8007C0078003E7C007F800F800F9FFCF3FBFF1F9FF9FF;
defparam sdpb_inst_5.INIT_RAM_02 = 256'h000003FFFFFF8000000000000000003FFFFFFFF9FF9F3FF9E003F3FFFE1FFE00;
defparam sdpb_inst_5.INIT_RAM_03 = 256'h078F000FE003E001E7FF1C7C7F87E7FC7FFFFFFFFFFFFFFFFFFFFFFFFFFE0000;
defparam sdpb_inst_5.INIT_RAM_04 = 256'h03FFFFFFFE3FE3CFFC7800FCFFFF87FF800FFC3FF800FFF8FF8FFC000E001E00;
defparam sdpb_inst_5.INIT_RAM_05 = 256'hFF9FFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000FFFFFFF80000000000000000;
defparam sdpb_inst_5.INIT_RAM_06 = 256'hFFC0E3FF07FE1C1FFF3FE3FFC007E003C003E3C00FF038FC4078FFCF1F1FE1F9;
defparam sdpb_inst_5.INIT_RAM_07 = 256'hF0000000003FFFFFFF8000000000000000007FFFFFFF8FF8F1FF1F003F1FFFE1;
defparam sdpb_inst_5.INIT_RAM_08 = 256'hF8FF8FF8F8FFFC7F3FFF1F3FF3E7E3F83E3FE7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_09 = 256'h0000000FFFFFFFF1FE3C7FC7FF87C7FFF83FF1FC7FC1FF8FC3FFC7FCFFFF1FFF;
defparam sdpb_inst_5.INIT_RAM_0A = 256'hFE0F8FF8FFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFFF00000000000;
defparam sdpb_inst_5.INIT_RAM_0B = 256'hFFFE0FF87F1FF07FE7F8FFF1FF1FFFE7FFFE3FE3FF3E3FFF3FC7FFE3C7FCF8F8;
defparam sdpb_inst_5.INIT_RAM_0C = 256'hFFFFFF0000000001FFFFFFFE000000000000000000FFFFFFFC7FC78FF1FFF1F1;
defparam sdpb_inst_5.INIT_RAM_0D = 256'hF8FFFF8FF8FFCFC7FFCFF1FFF8F1FF3E3F3F83E3FE3FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0E = 256'h0000000000001FFFFFFF1FF1E3FC7FFC7C3FFF81FF1FC7FC0FF9FE3FFE7FC7FF;
defparam sdpb_inst_5.INIT_RAM_0F = 256'hCF8FCFE4FC7F8FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFE00000;
defparam sdpb_inst_5.INIT_RAM_10 = 256'hFF9F8FFFE27FC7F9FF03FF7FC7FF9FF9FFFE3FFFE1FF1FF1F8FFF3FC7FFE3E3F;
defparam sdpb_inst_5.INIT_RAM_11 = 256'hFFFFFFFFFFF8000000000FFFFFFFFC000000000000000003FFFFFFC7FC7CFF1F;
defparam sdpb_inst_5.INIT_RAM_12 = 256'hFE7FFF8FFFFC7FC7FC7E3FFC7F8FFF8F8FF3E3F3F93F1FF1FFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_13 = 256'h0000000000000000007FFFFFF9FF9F1FC7FFE3E3FFF99FF1FE7FC67FFFF1FFE7;
defparam sdpb_inst_5.INIT_RAM_14 = 256'hF3F3FCFCFCFE4FC7FC7FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000003FFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_15 = 256'hE7F1FFF8FCFFFE63FE7F8FF19FFFFC7FF8FF9FFFF3FFFF1FF1FF1FC7FF1FE3FF;
defparam sdpb_inst_5.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFC000000000FFFFFFFFF000000000000000000FFFFFFE7FE7;
defparam sdpb_inst_5.INIT_RAM_17 = 256'h1FFE3FE3FFFCFFFFC7FE7FE7F0FFE3FCFFFC7C7F3F1F3F11F9FF1FFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_18 = 256'hFFFFFC000000000000000001FFFFFF8FF9F8FC7FFE3F3FFF9CFF9FE3FC67FFFF;
defparam sdpb_inst_5.INIT_RAM_19 = 256'hFF3FFF1F1FCFC7C7C47E7FE7FFFFFFFFFFFFFFFFFFFFFFFFFFF0000000003FFF;
defparam sdpb_inst_5.INIT_RAM_1A = 256'hE3FE3E3F1FFF8FCFFFE71FE7F8FF18FFFFC7FF8FF8FFFF1FFFF9FF9FF9FE3FF8;
defparam sdpb_inst_5.INIT_RAM_1B = 256'hE00000000000000007FFFE0000000007FFFFFFFF8000000000000000003FFFFF;
defparam sdpb_inst_5.INIT_RAM_1C = 256'h3FFFE1FFF1FE3FFFC7FFFC7FE7FE3FC7FF1FCFFF87E3F3F9F9F19F9FF9FFFFFF;
defparam sdpb_inst_5.INIT_RAM_1D = 256'h01FFFFFFFFF0000000000000000007FFFFFCFF8FC7C7FFE1F3FFF9E7F87E1FC7;
defparam sdpb_inst_5.INIT_RAM_1E = 256'hF1FFE3F3FFE1FCFC7E7E3C63E3FE7FFFFFF80000000000000000FFFF80000000;
defparam sdpb_inst_5.INIT_RAM_1F = 256'hFFFFFF3FF3F9F9FFF87C7FFE78FF8F87F1E7FFF0FFFC7FC7FFF1FFFF0FF8FF8F;
defparam sdpb_inst_5.INIT_RAM_20 = 256'hFFFFFE00000000000000001FFFE0000000003FFFFFFFFC000000000000000000;
defparam sdpb_inst_5.INIT_RAM_21 = 256'hE1FC79FFF03FFF1FF1FFFC7FF843FE3FE3FE3FF8787F007F3F1F9F8F38F8FF8F;
defparam sdpb_inst_5.INIT_RAM_22 = 256'h0000000FFFFFFFFF8000000000000000001FFFFFC7FCFE7E7F861F1FFF9F3FE1;
defparam sdpb_inst_5.INIT_RAM_23 = 256'h8FFCFFC7FF001FC00FC7C7E7F38F3E3FE3FFFFFFC00000000000000003FFF800;
defparam sdpb_inst_5.INIT_RAM_24 = 256'h000007FFFFF1FF1F8F9FE187E3FFE7CFFC007F1E3FF01FFFE7FC7FFF8FFE10FF;
defparam sdpb_inst_5.INIT_RAM_25 = 256'hC7F8FFFFFFF000000000000000007FFF0000000003FFFFFFFFF0000000000000;
defparam sdpb_inst_5.INIT_RAM_26 = 256'hF9FF001FC7CFF81FFFF9FF9FFFE3FF861FF1FF1FF1FFC007F063F8F1F8FCE3CF;
defparam sdpb_inst_5.INIT_RAM_27 = 256'hFFC0000000007FFFFFFFFC000000000000000000FFFFFC7FC7F1E7F801F8FFF9;
defparam sdpb_inst_5.INIT_RAM_28 = 256'hFF87FC7FC7FE3FF000FFF8FE3C7E3F38F3F1FF1FFFFFFE00000000000000001F;
defparam sdpb_inst_5.INIT_RAM_29 = 256'h00000000001FFFFF1FF1FC71FFFE7E3FFE3C3FC007F1F1FE0FFFFE7FE7FFFCFF;
defparam sdpb_inst_5.INIT_RAM_2A = 256'hCE7CFC7FC7FFFFFFFFFFFFFC0000000003FFF8000000001FFFFFFFFF80000000;
defparam sdpb_inst_5.INIT_RAM_2B = 256'h8FFF870FE1F9FC207F0FFFFF9FF9FFFF3FFFF1FF1FF9FF87F87E3FFE3FCF1F87;
defparam sdpb_inst_5.INIT_RAM_2C = 256'h0000FFFE0000000007FFFFFFFFE0000000000000000003FFFFE3FE7F9C7FFF8F;
defparam sdpb_inst_5.INIT_RAM_2D = 256'hFFCFFFFC7FE7FE7FF1FE3F8FFFC7F1C7F1F19F1F1FF1FFFFFFFFFFFFFF800000;
defparam sdpb_inst_5.INIT_RAM_2E = 256'h0000000000000000FFFFF8FF8FE71FFFE3F3FFE003F8FE3F000FC7FFFFE3FE7F;
defparam sdpb_inst_5.INIT_RAM_2F = 256'h71FC7C67C7E7FE7FFFFFFFFFFFFFF0000000001FFF8000000000FFFFFFFFF800;
defparam sdpb_inst_5.INIT_RAM_30 = 256'hFFF8FCFFF8007E3F8FC003F1FFFFF8FF8FFFF3FFFF9FF9FF9FFE3F8FF3FFF1FE;
defparam sdpb_inst_5.INIT_RAM_31 = 256'h0000000007FFE0000000003FFFFFFFFF0000000000000000001FFFFE3FE3F8C7;
defparam sdpb_inst_5.INIT_RAM_32 = 256'h1FE3FFFC7FFFE7FE7FE7FF87E3FCFFFC7F8C7F9F99F8F9FF9FFFFFFFFFFFFFFE;
defparam sdpb_inst_5.INIT_RAM_33 = 256'hFFC0000000000000000007FFFFCFF8FF19FFFE1F1FFE3F0F8FF1F0F8FC7FFFFF;
defparam sdpb_inst_5.INIT_RAM_34 = 256'hFF9FE31FE7E27E3E3FE7FFFFFFFFFFFFFFC000000001FFFC000000000FFFFFFF;
defparam sdpb_inst_5.INIT_RAM_35 = 256'h3FC47FFFC7C7EF8FE3F3FC7C7F1F1FFFFFC7FCFFFF1FFFF8FF8FF8FFF1F8FF3F;
defparam sdpb_inst_5.INIT_RAM_36 = 256'hFFFFF8000000003FFF0000000001FFFFFFFFF0000000000000000000FFFFF3FF;
defparam sdpb_inst_5.INIT_RAM_37 = 256'hFE7FF1FF1FFFC3FFFE3FE3FE3FFE3E3FC7FFE7FC07F9F89F8F8FF8FFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_38 = 256'hFFFFFFFE0000000000000000001FFFFCFFCFF81FFFF1F1F9E3FCFCFF1F1FE3C7;
defparam sdpb_inst_5.INIT_RAM_39 = 256'hC7F1FFF9FF81FE7E07F3F3FE3FFFFFFFFFFFFFFF000000000FFFE0000000007F;
defparam sdpb_inst_5.INIT_RAM_3A = 256'hFF1FF3FE07FFFC7E7E38FF1F3FC7C7F8F1FF1FFC7FC7FFF8FFFF8FF8FFC7FF8F;
defparam sdpb_inst_5.INIT_RAM_3B = 256'hFFFFFFFFFFC000000001FFF8000000001FFFFFFFFF80000000000000000007FF;
defparam sdpb_inst_5.INIT_RAM_3C = 256'hFF3E7FC7FF9FF1FFFE3FFFE1FF1FF1FFF1F1FE7FFE3FE07F8F81FCFC7F8FFFFF;
defparam sdpb_inst_5.INIT_RAM_3D = 256'h0003FFFFFFFFE0000000000000000000FFFFC7FCFFC1FFFF9F8F8E7FC7CFF9F1;
defparam sdpb_inst_5.INIT_RAM_3E = 256'h7FFC3C7F9FFF8FF81FE3F07F3F0FE3FFFFFFFFFFFFFFF8000000007FFE000000;
defparam sdpb_inst_5.INIT_RAM_3F = 256'h001FFFF8FF3FF07FFFE7E3E39FF9F1FE7C7FC78FF1FFE3FC7FFF8FFFFC7FC7FC;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_21}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b0;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFF000000001FFFC000000000FFFFFFFFF80000000000000000;
defparam sdpb_inst_6.INIT_RAM_01 = 256'h7F8F1FF9F1F87FFC7E1FFFF3FFFF1FF1FF9FFF8F1FE3FFE1FF07FC7C3FC7E3F8;
defparam sdpb_inst_6.INIT_RAM_02 = 256'h000000001FFFFFFFFE00000000000000000007FFFF1F8FFE1FFFF8FC78E7FE3C;
defparam sdpb_inst_6.INIT_RAM_03 = 256'hFE7FE7FFC3E7F8FFF87FC3FF1F0FF1F87C3FFFFFFFFFFFFFFFC000000007FFF0;
defparam sdpb_inst_6.INIT_RAM_04 = 256'h00000001FFFFC7E3FF87FFFC3F1C39FFCF1FE3C7FE7C7E1FFF0F87FFFCFFFFC7;
defparam sdpb_inst_6.INIT_RAM_05 = 256'h7F001FFFFFFFFFFFFFFFF000000000FFFC0000000007FFFFFFFF800000000000;
defparam sdpb_inst_6.INIT_RAM_06 = 256'h7FF1C7F8F1FFDF800FFFE003FFFF3FF001FF9FF9F000F9FE3F001FF8FFC7E3FE;
defparam sdpb_inst_6.INIT_RAM_07 = 256'h3FFF8000000001FFFFFFFFF00000000000000000003FFFF800FFF1FF800FE01E;
defparam sdpb_inst_6.INIT_RAM_08 = 256'hFC007FE7FE7C001E7FCF8007FE3FF9F9FF9FF00FFFFFFFFFFFFFFFFE00000000;
defparam sdpb_inst_6.INIT_RAM_09 = 256'h00000000000007FFFF007FFC7FC003FC079FFE79FF3CFFF7F007FFFE01FFFFCF;
defparam sdpb_inst_6.INIT_RAM_0A = 256'hFF7FF7FE03FFFFFFFFFFFFFFFFC000000007FFE0000000007FFFFFFFFC000000;
defparam sdpb_inst_6.INIT_RAM_0B = 256'hFF03F7FFDEFFEFFFFFFE03FFFF807FFFFFFF003FFBFFFF000FBFF7F003FFDFFE;
defparam sdpb_inst_6.INIT_RAM_0C = 256'h000001FFFC000000000FFFFFFFFF00000000000000000001FFFFE03FFFBFF800;
defparam sdpb_inst_6.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000;
defparam sdpb_inst_6.INIT_RAM_0E = 256'h0000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFF0000000003FFFFFFFFC0;
defparam sdpb_inst_6.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_11 = 256'hFF800000000FFFC0000000007FFFFFFFF00000000000000000000FFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_13 = 256'hFFF800000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFF0000000001FFFFF;
defparam sdpb_inst_6.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_16 = 256'hFFFFFFFC00000000FFFE0000000007FFFFFFFE000000000000000000007FFFFF;
defparam sdpb_inst_6.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_18 = 256'hFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFF8000000000;
defparam sdpb_inst_6.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1B = 256'hFFFFFFFFFFFFE000000007FFF0000000003FFFFFFFE000000000000000000003;
defparam sdpb_inst_6.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1D = 256'h00000FFFFFFFF800000000000000000000FFFFFFFFFFFFFFFFDFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000001FFFC0000;
defparam sdpb_inst_6.INIT_RAM_1F = 256'h00003FFFFFFFFFFFFFFCE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFE000000003FFF0000000001FFFFFFFE0000000000000000;
defparam sdpb_inst_6.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_22 = 256'hE0000000007FFFFFFF800000000000000000000FFFFFFFFFFFFFFF11FFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000FFF;
defparam sdpb_inst_6.INIT_RAM_24 = 256'h0000000001FFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFF000000003FFF8000000000FFFFFFFE00000000000;
defparam sdpb_inst_6.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_27 = 256'h007FFE0000000003FFFFFFF0000000000000000000007FFFFFFFFFFFFFF81FFF;
defparam sdpb_inst_6.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000;
defparam sdpb_inst_6.INIT_RAM_29 = 256'h000000000000000FFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000001FFFC000000000FFFFFFFC000000;
defparam sdpb_inst_6.INIT_RAM_2B = 256'hC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2C = 256'h00000003FFF0000000003FFFFFFE0000000000000000000003FFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sdpb_inst_6.INIT_RAM_2E = 256'h00000000000000000000FFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFC0000000007FFFFFF80;
defparam sdpb_inst_6.INIT_RAM_30 = 256'hFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_31 = 256'hFFFF000000003FFF8000000001FFFFFFE0000000000000000000003FFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_32 = 256'hFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_33 = 256'hFFF80000000000000000000007FFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_34 = 256'hFEFFFC007FFFFE7FFE003FFFFFFFFFFFFFFFFFC00000000FFFE0000000003FFF;
defparam sdpb_inst_6.INIT_RAM_35 = 256'hFFE3FCFFFF80FFFFCFF8FFFCFF8FFF8007FF8001FFFE03FFFFE007FFC001FFF7;
defparam sdpb_inst_6.INIT_RAM_36 = 256'hFFFFFFFFF000000001FFF8000000000FFFFFFC0000000000000000000001FFE7;
defparam sdpb_inst_6.INIT_RAM_37 = 256'hC000FFE0003FFE003FFFE000FFE0003FF07E1FFE000FFFFF8FFF0003FFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_38 = 256'h03FFFFFE00000000000000000000003FF0FFF07E1FFF800FFFE1FC1FFE1FE3FF;
defparam sdpb_inst_6.INIT_RAM_39 = 256'h0FFC1F83FF8001FFFFC3FFC000FFFFFFFFFFFFFFFFFE000000007FFF00000000;
defparam sdpb_inst_6.INIT_RAM_3A = 256'h0FFC3FFC1F87FFE001FFF87E07FF87F07FF0003FF0000FFF8007FFF0003FF800;
defparam sdpb_inst_6.INIT_RAM_3B = 256'hFFFFFFFFFFFFFF800000000FFFC0000000007FFFFF8000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3C = 256'hFC1FFC000FFE0003FFC000FFFC000FFE0003FF83E0FFE0007FFFF0FFF0003FFF;
defparam sdpb_inst_6.INIT_RAM_3D = 256'h0000001FFFFFC00000000000000000000003FF0FFF83E1FFF0003FFE1F81FFE0;
defparam sdpb_inst_6.INIT_RAM_3E = 256'hFF8000FFF0783FF8001FFFFC1FFC000FFFFFFFFFFFFFFFFFE000000003FFF800;
defparam sdpb_inst_6.INIT_RAM_3F = 256'h000000FFC1FFE0787FFC0007FF83E07FF83F87FF8003FF8000FFF0003FFF0001;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_22}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b0;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'h03FFFFFFFFFFFFFFFFF800000000FFFE0000000007FFFFF00000000000000000;
defparam sdpb_inst_7.INIT_RAM_01 = 256'h1FFE0FE1FFF0007FF0003FFC0E07FFC0007FF0007FFC0F0FFF0007FFFF07FF80;
defparam sdpb_inst_7.INIT_RAM_02 = 256'hFF8000000000FFFFF000000000000000000000003FF07FFC0E1FFE0381FFE0F8;
defparam sdpb_inst_7.INIT_RAM_03 = 256'hF07C1FFFC0FFFF81C3FFFFC1FFFFE1FFFFF0FFFFFFFFFFFFFFFFFF000000001F;
defparam sdpb_inst_7.INIT_RAM_04 = 256'h000000000007FC1FFF8183FF81E07FF83E07FFC3F87FFFFC1FFFC0FFFE07C0FF;
defparam sdpb_inst_7.INIT_RAM_05 = 256'h7FFFFC3FFFFFFFFFFFFFFFFFC000000007FFE0000000003FFFFC000000000000;
defparam sdpb_inst_7.INIT_RAM_06 = 256'hFF0F80FFF0FE0FFFFF07FFF87FFF83F83FFC3F87FFF87FFFF070FFFFF83FFFF8;
defparam sdpb_inst_7.INIT_RAM_07 = 256'h0000FFFC0000000007FFFE000000000000000000000001FF87FFF060FFE0FE0F;
defparam sdpb_inst_7.INIT_RAM_08 = 256'hFF0FFF0FE1FFFE1FFFFE0C3FFFFE0FFFFE1FFFFF07FFFFFFFFFFFFFFFFF80000;
defparam sdpb_inst_7.INIT_RAM_09 = 256'h00000000000000007FE1FFFE083FF87F83FFC3C03FFC3F83FFFFE1FFFE1FFFE0;
defparam sdpb_inst_7.INIT_RAM_0A = 256'hFFFF87FFFFC1FFFFFFFFFFFFFFFFFE000000003FFF0000000001FFFF00000000;
defparam sdpb_inst_7.INIT_RAM_0B = 256'h1FF07FF0F00FFF0FE0FFFFF87FFF87FFF83FC3FFC3F83FFF87FFFF810FFFFF83;
defparam sdpb_inst_7.INIT_RAM_0C = 256'h800000000FFFE0000000007FFF8000000000000000000000000FF87FFF800FFF;
defparam sdpb_inst_7.INIT_RAM_0D = 256'hFFFE1FF07FF07E0FFFE0FFFFF003FFFFE0FFFFE0FFFFF07FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0E = 256'h0000000000000000000003FE1FFFF003FFFFFC1FFC3803FFC1F03FFFFE1FFFE1;
defparam sdpb_inst_7.INIT_RAM_0F = 256'hFCF03FFFF83FFFFC1FFFFFFFFFFFFFFFFFE000000003FFF8000000001FFFC000;
defparam sdpb_inst_7.INIT_RAM_10 = 256'h00FFFFFF87FF0E00FFF0000FFFFF03FFF87FFF87FE1FFC1F83FFF83FFFFE00FF;
defparam sdpb_inst_7.INIT_RAM_11 = 256'hFFFFFC000000007FFE0000000003FF80000000000000000000000000FF87FFFE;
defparam sdpb_inst_7.INIT_RAM_12 = 256'hFFFE1FFFE1FF87FF8000FFFE0FFFFF803FFE000FFFFE0FFF0007FFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_13 = 256'h800000000000000000000000003FE1FFFF801FFFFFE1FFC3803FFC0003FFE000;
defparam sdpb_inst_7.INIT_RAM_14 = 256'hE00FFF8003FFFFC3FFC001FFFFFFFFFFFFFFFFFF000000001FFFC0000000007F;
defparam sdpb_inst_7.INIT_RAM_15 = 256'h7FFFE007FFFFF87FF0E10FFF0000FFF0003FFF83FFF87FE0FFE0003FFFC3FFFF;
defparam sdpb_inst_7.INIT_RAM_16 = 256'hFFFFFFFFFFC000000003FFF000000000000000000000000000000000000007F8;
defparam sdpb_inst_7.INIT_RAM_17 = 256'hFE000FFFE0FFFE1FF83FFC000FFFF0FFFFF801FFE000FFFFF0FFF0003FFFFFFF;
defparam sdpb_inst_7.INIT_RAM_18 = 256'h00000000000000000000000000000001FE0FFFF001FFFFFE1FFC1843FFC0003F;
defparam sdpb_inst_7.INIT_RAM_19 = 256'h3FFFFC007FFC003FFFFC3FFC000FFFFFFFFFFFFFFFFFF800000000FFFC000000;
defparam sdpb_inst_7.INIT_RAM_1A = 256'h007F83FFFC007FFFFF87FF0430FFF0000FFF8003FFFC3FFF83FF0FFF0003FFFC;
defparam sdpb_inst_7.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFE000000003FFF800000000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_1C = 256'h0003FFF000FFFF0FFFE0FFC3FFC000FFFF0FFFFF001FFF000FFFFF0FFFC003FF;
defparam sdpb_inst_7.INIT_RAM_1D = 256'h0000000000000000000000000000000000001FF0FFFF001FFFFFE1FFE00C1FFC;
defparam sdpb_inst_7.INIT_RAM_1E = 256'h3FFFC3FFFF8007FFFFC1FFFFC3FFFFE0FFFFFFFFFFFFFFFFFFC000000007FFE0;
defparam sdpb_inst_7.INIT_RAM_1F = 256'h00000007FC3FFFC007FFFFF83FF80387FF03F0FFFFFC3FFFC3FFFC3FF0FFF000;
defparam sdpb_inst_7.INIT_RAM_20 = 256'hFC3FFFFFFFFFFFFFFFFFF000000001FFFC000000000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_21 = 256'hE1FFE0FC1FFFFF0FFFF07FFF0FFC3FFC1E0FFFF0FFFFE041FFFFF07FFFF0FFFF;
defparam sdpb_inst_7.INIT_RAM_22 = 256'h7FFF00000000000000000000000000000000000001FF0FFFE0C1FFFFFE0FFE00;
defparam sdpb_inst_7.INIT_RAM_23 = 256'hFF07C3FFFC1FFFF8387FFFFE1FFFFC3FFFFF0FFFFFFFFFFFFFFFFFFC00000000;
defparam sdpb_inst_7.INIT_RAM_24 = 256'h0000000000007FC3FFF8387FF8FF83FF80787FF87F87FFFFC3FFFC1FFFC3FF0F;
defparam sdpb_inst_7.INIT_RAM_25 = 256'h0FFFFFC3FFFFFFFFFFFFFFFFFF800000000FFFC0000000000000000000000000;
defparam sdpb_inst_7.INIT_RAM_26 = 256'hFFE01E1FFE1FE1FFFFF0FFFF07FFF07F83FFC3F07FFF87FFFE1E0FFFFF87FFFF;
defparam sdpb_inst_7.INIT_RAM_27 = 256'h000003FFF00000000000000000000000000000000000001FF07FFC0E1FFE1FE0;
defparam sdpb_inst_7.INIT_RAM_28 = 256'h1FE0FFF0FC1FFFE1FFFF0783FFFFE1FFFFC1FFFFF0FFFFFFFFFFFFFFFFFFE000;
defparam sdpb_inst_7.INIT_RAM_29 = 256'h000000000000000007FC1FFF0787FF83F83FF80787FF83F87FFFFC3FFFE1FFFC;
defparam sdpb_inst_7.INIT_RAM_2A = 256'h7FFFF07FFFFC3FFFFFFFFFFFFFFFFFFC000000007FFE0000000003FFFFFFE000;
defparam sdpb_inst_7.INIT_RAM_2B = 256'hE0FC1FFF03E0FFE0FE1FFFFF07FFF87FFF83F83FFC3F07FFF87FFFC1F0FFFFF8;
defparam sdpb_inst_7.INIT_RAM_2C = 256'hFF000000001FFF8000000000FFFFFFFE00000000000000000001FF87FFC1E1FF;
defparam sdpb_inst_7.INIT_RAM_2D = 256'h1FFFE07C0FFF0FE1FFFE1FFFE07C3FFC001FFF0C1FFF8E0FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2E = 256'hFFF00000000000000000007FE1FFE0783FF81E07FFC0F83FFC3F83FFC8C1FFFE;
defparam sdpb_inst_7.INIT_RAM_2F = 256'hFE0003FF0007FF0003FFFFFFFFFFFFFFFFFFC000000007FFF0000000003FFFFF;
defparam sdpb_inst_7.INIT_RAM_30 = 256'h3E0FFF0001FFF03E0FFF0FE0FFE0007FFF87FFFC0007FFC1F87FFF87FFF83F0F;
defparam sdpb_inst_7.INIT_RAM_31 = 256'hFFFFFFF000000001FFFC0000000007FFFFFFFE0000000000000000001FF87FF8;
defparam sdpb_inst_7.INIT_RAM_32 = 256'h1FFFE1FFFF0001FFF07E1FFFE1FFFE0FC3FF8000FFC001FFC0007FFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_33 = 256'hFFFFFFFFC0000000000000000007FE1FFE0FC3FFC0007FFC0FC3FFC3F83FF800;
defparam sdpb_inst_7.INIT_RAM_34 = 256'h07F0FFE0003FF0003FF0001FFFFFFFFFFFFFFFFFFE000000003FFF0000000001;
defparam sdpb_inst_7.INIT_RAM_35 = 256'h87FF03F0FFF8003FFF03F0FFF0FF0FFE0007FFF87FFFE000FFFC1F87FFF83FFF;
defparam sdpb_inst_7.INIT_RAM_36 = 256'hFFFFFFFFFFFF800000000FFFE0000000007FFFFFFFFC000000000000000001FF;
defparam sdpb_inst_7.INIT_RAM_37 = 256'hFF8000FFFE1FFFFC003FFF07E1FFFE0FFFC1FC3FF8000FFC000FFC0007FFFFFF;
defparam sdpb_inst_7.INIT_RAM_38 = 256'h00000FFFFFFFFF0000000000000000007FE1FFC1FC3FFF001FFFC1FC3FFC3FC3;
defparam sdpb_inst_7.INIT_RAM_39 = 256'hC3FFF07F0FFE0003FF0007FF8001FFFFFFFFFFFFFFFFFFF000000001FFF80000;
defparam sdpb_inst_7.INIT_RAM_3A = 256'h001FF87FF07F0FFFE007FFF07F0FFF0FF0FFE0007FFF87FFFF801FFFC1FC7FFF;
defparam sdpb_inst_7.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFC000000007FFE0000000003FFFFFFFFE000000000000000;
defparam sdpb_inst_7.INIT_RAM_3C = 256'hE7FE7FFC003FFFF3FFFFF00FFFF9FF1FFFFBFFFE3FF7FFC001FFF003FFF001FF;
defparam sdpb_inst_7.INIT_RAM_3D = 256'hC000000000FFFFFFFFFC000000000000000007FF3FFE3FE7FFFC03FFFE7FE7FF;
defparam sdpb_inst_7.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFF;
defparam sdpb_inst_7.INIT_RAM_3F = 256'h00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[30:0],sdpb_inst_8_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_23}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_8.READ_MODE = 1'b0;
defparam sdpb_inst_8.BIT_WIDTH_0 = 1;
defparam sdpb_inst_8.BIT_WIDTH_1 = 1;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_8.RESET_MODE = "SYNC";
defparam sdpb_inst_8.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFE000000003FFF0000000001FFFFFFFFF8000000000;
defparam sdpb_inst_8.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_02 = 256'h00FFFC0000000007FFFFFFFFF000000000000000007FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000;
defparam sdpb_inst_8.INIT_RAM_04 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFF8000000000FFFFFFFFFE0000;
defparam sdpb_inst_8.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_07 = 256'h00000007FFE0000000003FFFFFFFFF800000000000000007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sdpb_inst_8.INIT_RAM_09 = 256'hF00000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFF8000000000FFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0C = 256'hFFFE000000003FFF0000000003FFFFFFFFFC00000000000000007FFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0E = 256'hFFFFFF80000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFC000000000FFFF;
defparam sdpb_inst_8.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_11 = 256'hFFFFFFFFE000000003FFF8000000001FFFFFFFFFE00000000000000007FFFFFF;
defparam sdpb_inst_8.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_13 = 256'h07FFFFFFFFF80000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFE00000000;
defparam sdpb_inst_8.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_16 = 256'hFFFFFFFFFFFFFF000000001FFF8000000001FFFFFFFFFF0000000000000000FF;
defparam sdpb_inst_8.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_18 = 256'h0000007FFFFFFFFFE0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000003FFF000;
defparam sdpb_inst_8.INIT_RAM_1A = 256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFF800000000FFFC000000000FFFFFFFFFF8000000000000;
defparam sdpb_inst_8.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1D = 256'hFF8000000003FFFFFFFFFE0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003F;
defparam sdpb_inst_8.INIT_RAM_1F = 256'h00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFE000000000FFFFFFFFFF80000000;
defparam sdpb_inst_8.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_22 = 256'h0001FFF8000000003FFFFFFFFFF0000000000000003FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000;
defparam sdpb_inst_8.INIT_RAM_24 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1FFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_25 = 256'hFFE1FF000FFFFFFFFFFFFFFFFFFFFC000000007FFE000000000FFFFFFFFFFC00;
defparam sdpb_inst_8.INIT_RAM_26 = 256'h3FC7FFFE1FFF8007FF07FFC01FFFFE3F87FFFC001F8007E0007FE3FC7F0F87F1;
defparam sdpb_inst_8.INIT_RAM_27 = 256'h000000001FFFC000000003FFFFFFFFFF0000000000000007FFFE3F8FC7FC7C00;
defparam sdpb_inst_8.INIT_RAM_28 = 256'h0FE1FFFE0003C001F0001FF87E1FC3E0F83FF03FC001FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_29 = 256'hFFC000000000000001FFFF0FE1F0FE1F0007E1FFFF03FFC001FFC1FFE003FFFF;
defparam sdpb_inst_8.INIT_RAM_2A = 256'hF81F0FFC0FF0007FFFFFFFFFFFFFFFFFFFE000000003FFF000000000FFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2B = 256'h87C001F87FFFC0FFF0007FE07FF8007FFFC1F87FFF8000F0003C0007FE1F83F0;
defparam sdpb_inst_8.INIT_RAM_2C = 256'hFFFFF800000000FFFE000000003FFFFFFFFFF0000000000000007FFFC1F87C1F;
defparam sdpb_inst_8.INIT_RAM_2D = 256'h1FFFF07E0FFFF0003E000F8001FF87F0FC3F03C3FF01FC001FFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2E = 256'hFFFFFFFC000000000000001FFFF07E0F07E1F0007E0FFFF01FF8001FF80FFE00;
defparam sdpb_inst_8.INIT_RAM_2F = 256'hFC3F0FE0F0FFC07F8007FFFFFFFFFFFFFFFFFFFF000000001FFF800000000FFF;
defparam sdpb_inst_8.INIT_RAM_30 = 256'h83E1F87C001FC3FFFC07FE0003FE03FF8383FFFE1FC3FFFC000F8003E0007FE0;
defparam sdpb_inst_8.INIT_RAM_31 = 256'hFFFFFFFFFFC000000007FFE000000003FFFFFFFFFF000000000000000FFFFE1F;
defparam sdpb_inst_8.INIT_RAM_32 = 256'h7FE1E0FFFF87F0FFFF0007E000FC001FFC3F0FC1FC1C3FF01FFFE1FFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_33 = 256'h00FFFFFFFFFFE000000000000003FFFF87F0F87E1F8003F0FFFF01FF8000FF80;
defparam sdpb_inst_8.INIT_RAM_34 = 256'h7FFF0FC3F87F8307FC03FFF83FFFFFFFFFFFFFFFFFFFF000000001FFFC000000;
defparam sdpb_inst_8.INIT_RAM_35 = 256'hFFE1FC3E0F87FFE0FC3FFFC03FE0F83FE01FF87C3FFFE1FC3FFFFE0FFFFC1FF0;
defparam sdpb_inst_8.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFC000000003FFF000000003FFFFFFFFFF800000000000000FF;
defparam sdpb_inst_8.INIT_RAM_37 = 256'h0FF807FE3F07FFF83F0FFFFF87FFFF87FE1FFFC3F0FE1FE0E1FF00FFFF0FFFFF;
defparam sdpb_inst_8.INIT_RAM_38 = 256'h0000000FFFFFFFFFFE000000000000003FFFF83F0FC3E1FFFC3F0FFFF00FF87F;
defparam sdpb_inst_8.INIT_RAM_39 = 256'hE1FF87FFF0FC3F87FC007FC03FFFC3FFFFFFFFFFFFFFFFFFFF800000000FFFC0;
defparam sdpb_inst_8.INIT_RAM_3A = 256'h001FFFFF0FC3F0787FFF0FC1FFFC21FE1FC3FE00FF8FC1FFFF0FC3FFFFE0FFFF;
defparam sdpb_inst_8.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFE000000001FFF800000003FFFFFFFFFF000000000000;
defparam sdpb_inst_8.INIT_RAM_3C = 256'h7F87F0FF803FFFE07FFFC3F0FFFFFC3FFFF87FE1FFFC3F0FE1FF801FF007FFF0;
defparam sdpb_inst_8.INIT_RAM_3D = 256'h7FFE00000000FFFFFFFFFFC000000000000007FFFFC3F0FE1E1FFFC3F87FFF08;
defparam sdpb_inst_8.INIT_RAM_3E = 256'h0FFFFC1FF87FFF0FC1F83FF007F861FFFC3FFFFFFFFFFFFFFFFFFFFC00000000;
defparam sdpb_inst_8.INIT_RAM_3F = 256'h00000001FFFFF0FC3F8787FFF07E1FFFC21FF0FC3FE187FFF81FFFF0FC1FFFFF;

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[30:0],sdpb_inst_9_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_9}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_24}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_9.READ_MODE = 1'b0;
defparam sdpb_inst_9.BIT_WIDTH_0 = 1;
defparam sdpb_inst_9.BIT_WIDTH_1 = 1;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_9.RESET_MODE = "SYNC";
defparam sdpb_inst_9.INIT_RAM_00 = 256'h3F800FFFFFFFFFFFFFFFFFFFFF000000001FFF800000003FFFFFFFFFF0000000;
defparam sdpb_inst_9.INIT_RAM_01 = 256'hFFF083FC1F07F861FFF007FFFC3F07FFFFC3FF8007FE1FFFC1F87F0FFC01FE18;
defparam sdpb_inst_9.INIT_RAM_02 = 256'h000007FFF00000000FFFFFFFFFFC00000000000000FFFFFC3F87E1E1FE001F87;
defparam sdpb_inst_9.INIT_RAM_03 = 256'hFFFFF0FFE001FF83FFF87E1FC3FF007F870FE001FFFFFFFFFFFFFFFFFFFFC000;
defparam sdpb_inst_9.INIT_RAM_04 = 256'h0000000000003FFFFF0FE1FC387F0007E1FFFC30FF8001FE187FF001FFFF0FE1;
defparam sdpb_inst_9.INIT_RAM_05 = 256'h1FE1C3F8007FFFFFFFFFFFFFFFFFFFF800000000FFFC00000007FFFFFFFFFF00;
defparam sdpb_inst_9.INIT_RAM_06 = 256'h01F87FFF0E1FE0007F860FF800FFFFC3F87FFFFC3FF8007FE0FFFE1F87F0FFC0;
defparam sdpb_inst_9.INIT_RAM_07 = 256'hFE000000003FFF00000001FFFFFFFFFFC00000000000000FFFFFC3F87F0E1FC0;
defparam sdpb_inst_9.INIT_RAM_08 = 256'hF0FE1FFFFF0FFE000FFC3FFF87E0FC3FF003F8787E001FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_09 = 256'hFFE000000000000007FFFFF0FE1FC387F0007E1FFFC387F8001FE1C3FC007FFF;
defparam sdpb_inst_9.INIT_RAM_0A = 256'h0FF800FE1E1F8007FFFFFFFFFFFFFFFFFFFF8000000007FFC00000007FFFFFFF;
defparam sdpb_inst_9.INIT_RAM_0B = 256'h61FE001F87FFF0E1FF0007F870FF003FFFFC1F83FFFFC3FFC003FF0FFFE1FC3F;
defparam sdpb_inst_9.INIT_RAM_0C = 256'hFFFFFFF000000001FFF00000003FFFFFFFFFF800000000000001FFFFFC3F83F8;
defparam sdpb_inst_9.INIT_RAM_0D = 256'h1FFFFF87F0FFFFF87FF800FFC3FFF87F0FC3FE003F8383F001FFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_0E = 256'hFFFFFFFE00000000000000FFFFFF07E0FE18FFC003E0FFFC387FC001FE1C1FC0;
defparam sdpb_inst_9.INIT_RAM_0F = 256'h1FC3F0FF820FE000FFF87FFFFFFFFFFFFFFFFFFFFC000000007FF80000000FFF;
defparam sdpb_inst_9.INIT_RAM_10 = 256'hFC3FC03FFFE0FC3F7F0C0FF0007F8007E01FFFFFE1FC3FFFFE1FFFFC3FF0FFFE;
defparam sdpb_inst_9.INIT_RAM_11 = 256'hFFFFFFFFFFFF000000000FFE00000003FFFFFFFFFF000000000000003FFFFFE1;
defparam sdpb_inst_9.INIT_RAM_12 = 256'h00F81FFFFFF87F0FFFFF87FFFF0FFC3FFF83F0FC3FC1C3F8003FFE1FFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_13 = 256'h00FFFFFFFFFFC00000000000001FFFFFF87F0FF00FFFFC3F0F1FC003F81E0FC0;
defparam sdpb_inst_9.INIT_RAM_14 = 256'h0FFFF0FC3F07F0707E000FFF87FFFFFFFFFFFFFFFFFFFFC000000001FF000000;
defparam sdpb_inst_9.INIT_RAM_15 = 256'hFFFE1FC3FC03FFFF0FC3C3F0007E0F83F0003F0FFFFFFE0FC3FFFFE1FFFFC3FF;
defparam sdpb_inst_9.INIT_RAM_16 = 256'hFFFFFFFFFE000000000000000000000000007FFFFFFFFFE000000000000007FF;
defparam sdpb_inst_9.INIT_RAM_17 = 256'hF0FC000FC3F87FFFC3F0FFFFF83FFFF0FFC1FFFC3F07C1FC1E1F8001FFF0FFFF;
defparam sdpb_inst_9.INIT_RAM_18 = 256'h0000003FFFFFFFFFF800000000000003FFFFFFC3F0FF80FFFFC3F0F0F8001F83;
defparam sdpb_inst_9.INIT_RAM_19 = 256'hFE1FF87FFF0FC1F07F0F87E0007FFC3FFFFFFFFFFFFF00000000000000000000;
defparam sdpb_inst_9.INIT_RAM_1A = 256'h00FFFFFFF0FC3FE03FFFF0FE1C3E0003F0FC3F0003F0FE1FFFF0FC3FFFFF0FFF;
defparam sdpb_inst_9.INIT_RAM_1B = 256'h0FFFFFFFFFFFFFC00000000000000000000000000FFFFFFFFFFC000000000000;
defparam sdpb_inst_9.INIT_RAM_1C = 256'h00FC3F0FC0007C1F07FFFC1F0FFFFFC3FFFF07FE1FFF83F83C1F83E1F8000FFF;
defparam sdpb_inst_9.INIT_RAM_1D = 256'h000000000007FFFFFFFFFE000000000000007FFFFFFC3F0FF80FFFFC3F870F80;
defparam sdpb_inst_9.INIT_RAM_1E = 256'hF0FFC001FF87F0007E0607E0F87E0F83FFC3FFFFFFFFFFFFF000000000000000;
defparam sdpb_inst_9.INIT_RAM_1F = 256'h0000003FFFFFFF0383FF03FF000FE0C1E0FC3F0FC1F07C0F8381FFFF0303FFFF;
defparam sdpb_inst_9.INIT_RAM_20 = 256'hF0FFF07FFFFFFFFFFFFC00000000000000000000000003FFFFFFFFFF80000000;
defparam sdpb_inst_9.INIT_RAM_21 = 256'h20787F0FC3F87C3FC3E0007FFFE000FFFFFC3FF0007FE1FC001FC001F83E1F87;
defparam sdpb_inst_9.INIT_RAM_22 = 256'h0000000000000001FFFFFFFFFF800000000000001FFFFFFFE000FFC0FF8001F8;
defparam sdpb_inst_9.INIT_RAM_23 = 256'h3FFFFF0FFC001FF83F0007F000FC1F87E1FC1FFE1FFFFFFFFFFFFF8000000000;
defparam sdpb_inst_9.INIT_RAM_24 = 256'h000000000007FFFFFFF8003FF03FE0007E003E1FE1F07E1F0FF0F8001FFFF800;
defparam sdpb_inst_9.INIT_RAM_25 = 256'hE1F87F87FF87FFFFFFFFFFFFFFFFFFFFE000000001FFFFFFFFFFFFFFFFFFC000;
defparam sdpb_inst_9.INIT_RAM_26 = 256'h001FC00F87F83C1F87C3FC3F000FFFFF001FFFFFC3FF0003FF0FC001FE003F07;
defparam sdpb_inst_9.INIT_RAM_27 = 256'hFFF800000000FFFFFFFFFFFFFFFFFFF000000000000003FFFFFFFF000FFE0FF8;
defparam sdpb_inst_9.INIT_RAM_28 = 256'hFFE007FFFFF0FFC000FFC3F0007FC00FC1FC7E1FE1FFE1FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_29 = 256'hF000000000000001FFFFFFFFC007FF83FE0007F803E1FF0F07E1F0FF07E007FF;
defparam sdpb_inst_9.INIT_RAM_2A = 256'h07F8FF1FCFFC7FFCFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2B = 256'hF1FFC003FE01F8FFC7E3FC7C7FE3FC01FFFFF803FFFFFE3FF0007FF1FE001FF8;
defparam sdpb_inst_9.INIT_RAM_2C = 256'hFFFFFFFFC000000003FFFFFFFFFFFFFFFFF000000000000001FFFFFFFFF803FF;
defparam sdpb_inst_9.INIT_RAM_2D = 256'hE3FFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2E = 256'hFFFFF8000000000000007FFFFFFFFFC3FFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFFFFFE000000001FFFFFFF8000000000000000000000007FFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_33 = 256'h0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000;
defparam sdpb_inst_9.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000001FFFFF;
defparam sdpb_inst_9.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_38 = 256'h00000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000;
defparam sdpb_inst_9.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000003F;
defparam sdpb_inst_9.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3D = 256'h000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000;
defparam sdpb_inst_9.INIT_RAM_3F = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_10 (
    .DO({sdpb_inst_10_dout_w[30:0],sdpb_inst_10_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_10}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_25}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_10.READ_MODE = 1'b0;
defparam sdpb_inst_10.BIT_WIDTH_0 = 1;
defparam sdpb_inst_10.BIT_WIDTH_1 = 1;
defparam sdpb_inst_10.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_10.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_10.RESET_MODE = "SYNC";
defparam sdpb_inst_10.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000;
defparam sdpb_inst_10.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_02 = 256'h000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_04 = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000;
defparam sdpb_inst_10.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_07 = 256'hFFFFF000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0C = 256'hFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000001FFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFF;
defparam sdpb_inst_10.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000;
defparam sdpb_inst_10.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1D = 256'h000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam sdpb_inst_10.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_22 = 256'hFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_27 = 256'hFFFFFFE000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2C = 256'hFFFFFFFFFFFE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFF;
defparam sdpb_inst_10.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_38 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000;
defparam sdpb_inst_10.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3D = 256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam sdpb_inst_10.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_11 (
    .DO({sdpb_inst_11_dout_w[30:0],sdpb_inst_11_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_11}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_26}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_11.READ_MODE = 1'b0;
defparam sdpb_inst_11.BIT_WIDTH_0 = 1;
defparam sdpb_inst_11.BIT_WIDTH_1 = 1;
defparam sdpb_inst_11.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_11.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_11.RESET_MODE = "SYNC";
defparam sdpb_inst_11.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_02 = 256'hFFF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_07 = 256'hFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000001FFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0C = 256'hFFFFFFFFFFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000FFFFFFF;
defparam sdpb_inst_11.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFE000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FF;
defparam sdpb_inst_11.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_18 = 256'h0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam sdpb_inst_11.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1D = 256'h000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_11.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_22 = 256'hFFFFE000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_27 = 256'hFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFF000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFFFF;
defparam sdpb_inst_11.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFF8000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001;
defparam sdpb_inst_11.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_38 = 256'h00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam sdpb_inst_11.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3D = 256'hF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_12 (
    .DO({sdpb_inst_12_dout_w[30:0],sdpb_inst_12_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_12}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_27}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_12.READ_MODE = 1'b0;
defparam sdpb_inst_12.BIT_WIDTH_0 = 1;
defparam sdpb_inst_12.BIT_WIDTH_1 = 1;
defparam sdpb_inst_12.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_12.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_12.RESET_MODE = "SYNC";
defparam sdpb_inst_12.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000001FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_02 = 256'hFFFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_07 = 256'hFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFE000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000007FFF;
defparam sdpb_inst_12.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_13 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000;
defparam sdpb_inst_12.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_18 = 256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam sdpb_inst_12.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1D = 256'hFFF000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_22 = 256'hFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_27 = 256'hFFFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000001FFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FF;
defparam sdpb_inst_12.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_33 = 256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000;
defparam sdpb_inst_12.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_38 = 256'h000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_12.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3D = 256'hFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_13 (
    .DO({sdpb_inst_13_dout_w[30:0],sdpb_inst_13_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_13}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_28}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_13.READ_MODE = 1'b0;
defparam sdpb_inst_13.BIT_WIDTH_0 = 1;
defparam sdpb_inst_13.BIT_WIDTH_1 = 1;
defparam sdpb_inst_13.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_13.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_13.RESET_MODE = "SYNC";
defparam sdpb_inst_13.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000FFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_02 = 256'hFFFFFFFFFE000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFF000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFFFF;
defparam sdpb_inst_13.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFF800000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003;
defparam sdpb_inst_13.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_13 = 256'h00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam sdpb_inst_13.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000007FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_18 = 256'hF800000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000003FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1D = 256'hFFFFFFC00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000003FFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_22 = 256'hFFFFFFFFFFFE000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000001FFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFF000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000FFFF;
defparam sdpb_inst_13.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFF800000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2E = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000;
defparam sdpb_inst_13.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_33 = 256'h0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam sdpb_inst_13.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_38 = 256'hFFF800000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3D = 256'hFFFFFFFFC00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_14 (
    .DO({sdpb_inst_14_dout_w[30:0],sdpb_inst_14_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_14}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_29}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_14.READ_MODE = 1'b0;
defparam sdpb_inst_14.BIT_WIDTH_0 = 1;
defparam sdpb_inst_14.BIT_WIDTH_1 = 1;
defparam sdpb_inst_14.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_14.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_14.RESET_MODE = "SYNC";
defparam sdpb_inst_14.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_02 = 256'hFFFFFFFFFFFFFF00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000003FFFFFFF;
defparam sdpb_inst_14.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFF80000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FF;
defparam sdpb_inst_14.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0E = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000;
defparam sdpb_inst_14.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_13 = 256'hC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000003FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_18 = 256'hFFFFFF00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000001FFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1D = 256'hFFFFFFFFFFFC0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000FFFFFF;
defparam sdpb_inst_14.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007;
defparam sdpb_inst_14.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2E = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sdpb_inst_14.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_33 = 256'hFFFFC00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_38 = 256'hFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3F = 256'h000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[17]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[16]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[15]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sdpb_inst_2_dout[0]),
  .I1(sdpb_inst_3_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sdpb_inst_4_dout[0]),
  .I1(sdpb_inst_5_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sdpb_inst_6_dout[0]),
  .I1(sdpb_inst_7_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(sdpb_inst_8_dout[0]),
  .I1(sdpb_inst_9_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(sdpb_inst_10_dout[0]),
  .I1(sdpb_inst_11_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sdpb_inst_12_dout[0]),
  .I1(sdpb_inst_13_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_2)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_2)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_2)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_6),
  .I1(sdpb_inst_14_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_1)
);
MUX2 mux_inst_14 (
  .O(dout[0]),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_0)
);
endmodule //Gowin_SDPB3
