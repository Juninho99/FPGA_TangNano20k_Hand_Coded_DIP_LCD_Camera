//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Wed Aug 23 13:45:11 2023

module Gowin_SDPB2 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);//gaussian_blur_5x5

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [13:0] ada;
input [7:0] din;
input [13:0] adb;

wire [29:0] sdpb_inst_0_dout_w;
wire [1:0] sdpb_inst_0_dout;
wire [29:0] sdpb_inst_1_dout_w;
wire [3:2] sdpb_inst_1_dout;
wire [29:0] sdpb_inst_2_dout_w;
wire [5:4] sdpb_inst_2_dout;
wire [29:0] sdpb_inst_3_dout_w;
wire [7:6] sdpb_inst_3_dout;
wire [23:0] sdpb_inst_4_dout_w;
wire [7:0] sdpb_inst_4_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[29:0],sdpb_inst_0_dout[1:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[13]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 2;
defparam sdpb_inst_0.BIT_WIDTH_1 = 2;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7D9FFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1BFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FF7FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFAFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFEEFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFC3FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCBFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF3FFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF9FFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFCFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFBFFEBFFFFA5FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFF8000000003FFF0000C3B2EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h34BE88FBF3FC000000003FFFEAA3FFFFE06BFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hB170CF6F3FEBFFFFFFFEFFF8004BFFFFFF3FFD83E823F7E0FFEFFB7D9432393B;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h3ABDB067FFFFFFFFFFFFFFEFFFBFFFFFFAFFCBEF6AFF2FEB7F2FF3DEA5B17710;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hDF94A3AFFEAAAA29EDFFFEFFFEFFFFFFCFFDF7BFEEF8ED7AEFF34FAFF9BBBB8F;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h6A673BFFEFFEFEB8EBFFEBFFFBFFFFFF9FDBB5E6BF8C07D60F3FFB93937DCDCA;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h2D23FFFFFFCFFFFFFFFF2FFFFFFFFFFEBFBA8F8AFEFC707DF3FFCEAAFB0CDED6;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h5F42FFFFFFBFFFFDFFFFFFFFFFFFFFFFFAEFFF1E3A7A227FCEFEFEB3FC2D3A8B;
defparam sdpb_inst_0.INIT_RAM_20 = 256'hFBEFFFFFFFFFEBC3FFFFFF7FFFFFFF7F86FF614B97FF4EFD6F8F1F73C856DB71;
defparam sdpb_inst_0.INIT_RAM_21 = 256'hFFFFFFFFDBFF7EFFFEBFFFFFFFFFFCFFEFAFAFFFEEBEBFFFFFEFFF6FFFFFFFFE;
defparam sdpb_inst_0.INIT_RAM_22 = 256'hFFFFFFFFBFFFF3FFCBFF3FFFFFFFCFFFFFF6FFFFFFFFFFEFFBFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_23 = 256'hFFFFFFFBFFCFBFFFFFDBFFFFFFFEFEFFFF4FFBFFFFFFEFFFFBFFFFFBFFBFFFBB;
defparam sdpb_inst_0.INIT_RAM_24 = 256'hFFFFFF7FFEEFFFFAEFBFFFFFFFFFE97FEDBE87F97C0D02C3BD0FD0823C3FCF81;
defparam sdpb_inst_0.INIT_RAM_25 = 256'hFFFFF9FFFFBFFF4F2FFFFFFFFFF3E4BEDFAFFD9730CCFEDB56B64C4731FC3FEF;
defparam sdpb_inst_0.INIT_RAM_26 = 256'hFFFFDFFF7EFFFFBABFFFFFFFFFEF33EEB84FC9FDCF1FF87FEFDFEC375FF7F7FF;
defparam sdpb_inst_0.INIT_RAM_27 = 256'hFFFDFFF7AFFFF0023FFFFFFF7EFFAFB3FFFCDBE0FBFBBEE9BD3EB384FF7F7FFF;
defparam sdpb_inst_0.INIT_RAM_28 = 256'hFFF7FFFFAFFF7FF4FFFFFFFBDF88CFBF77FEFE8F9FCF2CCBFFF13EDFF7FF3FFF;
defparam sdpb_inst_0.INIT_RAM_29 = 256'hFE7FFDEBFFFAFFF7FFFFFF7DF68E53C39B23C4FE7DC3CABF3EB7D8F5ED4BFFFF;
defparam sdpb_inst_0.INIT_RAM_2A = 256'hF3FFDF9FFFAFFFBFFFFFF3FF31FBFFAF97FFFFDFF82F93EBD27DF73FEFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2B = 256'hEFFC7EFFFAFFFDFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2C = 256'hFFFFEFFFDFFFFBFFFFF7FAEFEBFFFABFEEFFBFBABEFEFAFEFFAAAFBFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2D = 256'hFFBF3FFEFFFFFFFFFFBFA425CF9F5A76F7D7FFFFF33F8DE7DA19EF57FFFFFFFC;
defparam sdpb_inst_0.INIT_RAM_2E = 256'hFDFFFFEFFFF7FFFFF7FFC35E72F5BCACF83F98FD70BEBE31569C7C3FFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2F = 256'hEFBFFAFFFF7FFFFFBF7C9584CF2EB7C2B9FFC7F29FF7EBF3EFD083FFFFFFFF3F;
defparam sdpb_inst_0.INIT_RAM_30 = 256'hA7FF7FFFAFFFFFAFFDFD0FEDBAA85E381FFF3FBE8FFE68AD7E547FFFFFFFFBFF;
defparam sdpb_inst_0.INIT_RAM_31 = 256'hAA97FFF2FFFFFAFF4DFAB8F7A48FEEDAFFD7FDFCFEA39EA5D2F7FFFFF696AFFF;
defparam sdpb_inst_0.INIT_RAM_32 = 256'hFFFFF8BFFFFCFFFD8D497E4AC7CDA6CFE1BFFF3F8C3FD9ECFB8FFFFF3AAFFFF6;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h2FFFAFFFE6BFFFDDF696D61CEEEEE4FED3FCAAB16847DFBF36FFFFFFFFDFFFFF;
defparam sdpb_inst_0.INIT_RAM_34 = 256'hAAF3C5567BFFFFFFFFFFFFF7FFEBFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFF4EA;
defparam sdpb_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFE7FFF;
defparam sdpb_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFF;
defparam sdpb_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFF;
defparam sdpb_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FF9FFFFFF;
defparam sdpb_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFCFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFEFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF3FFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFEFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFF7FFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFEFFFFFFFFFFF;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[29:0],sdpb_inst_1_dout[3:2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[13]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 2;
defparam sdpb_inst_1.BIT_WIDTH_1 = 2;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE333FFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3F1BFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF7FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFF3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFEFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFDFFF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFC000000007FFFC000D3F1EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h305F6DEDFFFCFFFFFFFFFFFFFFFFFFFFF1BFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h5BFECC5F3FC555555556FFFD558FFFFFFF7FFFEFE837F3F0F7CBFBBC0C301C1E;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h7330D7FBFFFFFFFFFFFFFFFFFFFFFFFFFEFFFDBC1E3F9E7FFEBFF7D09E02A7DD;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hFBA6F37FFEAAAAEAFFFFFDFFFFFFFFFFCFFDD2DF9BF8EEF1FDF77FFFFCF2BCEF;
defparam sdpb_inst_1.INIT_RAM_1D = 256'hB7C33FFFFFFEFFFDFBFFFFFFFFFFFFFFFFCFE2CECFAEF3BFCF7EFFECFF7FF2FB;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h3A27CFFFFFF3FFFF3FFFBFFFFFFFFFFFFF7F6DFFFABDBC8BFDEFEDCEFBDC2FED;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h8EB4FFFFFFBFFFFCFFFBFFF3FFFFFFFFFFF6FCDCBB37F5BBCFFDFDF3BD9DBCCB;
defparam sdpb_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFF93FFFFFF7FFFFFFFFF73EF6913E7FFFB7FFFDF8F7B6BF14FB3;
defparam sdpb_inst_1.INIT_RAM_21 = 256'hFFFFFFFFEFFF7FFFFCFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFF7FFCFFFFFFFFFFFCFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_23 = 256'hFFFFFFF7FFCF3FFFBFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_24 = 256'hFFFFFF3FFDF7FFF3FFFFFFFFFFFF5DB3EFFCDBFCFC2C0BC9FE0FC3F9F80FEFC2;
defparam sdpb_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFBFFFFFF3FFFFFFFFF39F2FC87CF3CCBA7E6BE2FCEF99ECFE6FF7EBF;
defparam sdpb_inst_1.INIT_RAM_26 = 256'hFFFFEFFF7EFFFF3FFFFFFFFFF39FF7CBFCF3FD3DCFEFFE7CFFCBFBBD4FFFD5FF;
defparam sdpb_inst_1.INIT_RAM_27 = 256'hFFFEFFFFEFFFFAA9FFFFFFFF38FCFFF3C7BF3FF3FCFEF3D83DFFE3E1FF3E3FFF;
defparam sdpb_inst_1.INIT_RAM_28 = 256'hFFFFFFFFBFFFBFFCFFFFFFF3EFD3F7FFB7DD3FFFFFCBFE4BD3F87FDFF7FFBFFF;
defparam sdpb_inst_1.INIT_RAM_29 = 256'hFF7FFDFFFFFFFFF7FFFFFF3FF42FB7C7FF63D3FCFD1FC57F7EF3D274FE2BFFFF;
defparam sdpb_inst_1.INIT_RAM_2A = 256'hFBFFFFCFFF3FFFFFFFFFF7CF7EFA7F73EF3C0FDFF2FDFBF7F77D0F83E0BFFFFF;
defparam sdpb_inst_1.INIT_RAM_2B = 256'hDFFCBEFFFFFFFEFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2C = 256'hFFFFFFFFDFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFBF73F23BFFEFABEFC3FEFFC4F3DCFBF7F3F333FFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2E = 256'hFEF7FFDFFFF3FFFFFFFBED44FFF7FA3CBAFFDDFE02BDCF7F600EF93FFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2F = 256'hEFBFFFFFFFFFFFFEFFBC35F36F23BBE389FFFBF4EEBBFFA7DEC3EBFFFFFFFFBF;
defparam sdpb_inst_1.INIT_RAM_30 = 256'hB3FF3FFFEFFFFFCFF8DC2E5DFC3E2FFFCFEEBF9E2BBF3D1D9CFE3FFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h557BFFFBFFFFF7FF0EFAF5D98531C8FFFF73FEFC33F13FDBFBF9FFFFFFA97FFF;
defparam sdpb_inst_1.INIT_RAM_32 = 256'hFFFFFF7FFFFEBFFC5FFEDD7D62EEEF7FC53FFC7FAD2F8CFECFEFFFFF8552FFF1;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h75553FFFFEBFFFC7FBE9CA3FBECF55FF0FFCFF7DFEC58CCE7CFFFFFFFFFFFF3F;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h000415557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD55;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFF500;
defparam sdpb_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFF;
defparam sdpb_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFF3FFFFF;
defparam sdpb_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFEFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFCFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFF7FFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFDFFFFFFFFFFF;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[29:0],sdpb_inst_2_dout[5:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[13]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 2;
defparam sdpb_inst_2.BIT_WIDTH_1 = 2;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFED7FFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEADFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAA9FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAA3FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCAAABFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2AABFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6AAA3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAABFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAA9FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAA7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAA7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFCAAA8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFAAA8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF2AAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF6AAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFEAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFDAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFEAAAEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_18 = 256'hFFFFFFFFFFFFD55555555EAAA155503F09FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_19 = 256'hFFFFFFFFFFFCAAAAAAAAAAAAAAAAAAAAAD3FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1A = 256'h05F5DC8F7FFAAAAAAAABAAABFFAAAAAAA8BFFFFFFFFFFFFFFFFBFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1B = 256'hFBBADEFBFFFFFFFFFFDAAA8FFF2AAAAAA9FFDCCCCF7FFF0F3D0FB7C4CF32C1E3;
defparam sdpb_inst_2.INIT_RAM_1C = 256'h777EB77FF3FFFFFF3FAAA8FFFDAAAAAAB7FCFECFE7FCFEF3EEF7FF7FCEF6BEEF;
defparam sdpb_inst_2.INIT_RAM_1D = 256'h7B0337FFC000AAABFEAAAFFFFAAAAAAAAFEFBCE1EFDFEB0F9F7FFDD2EFBBEBCF;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h71FFEFFFFFFEAAAFAAAAFFFF2AAAAAABFFB74FBEFCF6F8E3FEFFDFAFBBEC8E8C;
defparam sdpb_inst_2.INIT_RAM_1F = 256'hFCC6FFFFFFAAAAFFAAAFFFF2AAAAAAAFFFFFFDEDEF77EAFBFFFEFCFF3E8FFDF7;
defparam sdpb_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFAAABDEAABFFF6AAAAAAABFDBCF59B3D3F379BF5FDF5B3E52FA6F3F;
defparam sdpb_inst_2.INIT_RAM_21 = 256'hFFFFFFFFDAAA7EAAA9FFFEAAAAAAA8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_22 = 256'hFFFFFFFFAAABFEAABFFF2AAAAAAA8FFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_23 = 256'hFFFFFFF6AAAFEAAABFFAAAAAAAAAFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_24 = 256'hFFFFFF6AABFEAAA3FCAAAAAAAAA77F33FBFCDFCCF43E03E9FC0FC3CEBC1FF7C0;
defparam sdpb_inst_2.INIT_RAM_25 = 256'hFFFFFEAAAFEAAABFAAAAAAAAAA31F2BEABCE7CDFBDEFFE7BFFFFFFAFF0FFBFEF;
defparam sdpb_inst_2.INIT_RAM_26 = 256'hFFFFDAAA3CAAA87AAAAAAAAAAFBFF3EFBDFBE2FE7FFFFFBFCFEBF6BEBFF3EBFF;
defparam sdpb_inst_2.INIT_RAM_27 = 256'hFFFEAAABFAAAA555EAAAAAAAFEFFBFF3E0FF97DBFFFFFFEFFD7F47EBFFFFBFFF;
defparam sdpb_inst_2.INIT_RAM_28 = 256'hFFFAAAAFEAAAFFFEAAAAAAAFCF9EF3FCFFDFFFEFEFCFBCC7F3FFFFDFFFFEFFFF;
defparam sdpb_inst_2.INIT_RAM_29 = 256'hFFEAAAFAAAABFFFEAAAAAAFEF24FDFFFBEF3F2FFFEDBEEFFBFBFC3F4BE37FFFF;
defparam sdpb_inst_2.INIT_RAM_2A = 256'hFEAAAFFAAAFFFFFAAAAAAFFFFFFDFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2B = 256'hFAAB7DAAABFFFDAAAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2C = 256'hAAA3FAAABFFFFAAAAAA3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2D = 256'hAABFEAAAFFFFAAAAAA3F7B7F977FDF97DFC7FDCFD5C4D1F73737DF47FFFFFFFC;
defparam sdpb_inst_2.INIT_RAM_2E = 256'hABFEAABFFFFEAAAAAFF3EB3EFAFEFAFFF9AFCFFE2EAEAFFB7ABDFFFFFFFFFFFA;
defparam sdpb_inst_2.INIT_RAM_2F = 256'hBFAAABFFFFAAAAABFFF9D3F39FD7FAFFF2FEFFF6FBFFFF31FDC7F3FFFFFFFF2A;
defparam sdpb_inst_2.INIT_RAM_30 = 256'h5AAA3FFFCAAAAA9FF6EC3C1FF7341F2CEFCFBFCE4BBFB3FD3F8C3FFFFFFFF6AA;
defparam sdpb_inst_2.INIT_RAM_31 = 256'h000FFFFEAAAAA7FFEFCBFDC61FAFF1FCFFE7FDFF76F2CDFCE2F6FFFFFD556AAA;
defparam sdpb_inst_2.INIT_RAM_32 = 256'hFFFFFCEAAAA9FFFF3FBD7FCBEDCCFF2FFD7FEF0BBC3EAFEFEBAFFFFFC003AAAC;
defparam sdpb_inst_2.INIT_RAM_33 = 256'h3FFFEAAAA83FFFFEF7D5FFBDDDEEF2FF8FFEF5BED6F3EEEFFEFFFFFFFFEAAAFF;
defparam sdpb_inst_2.INIT_RAM_34 = 256'hAAAAAAABBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAA800;
defparam sdpb_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAA;
defparam sdpb_inst_2.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAFFFF;
defparam sdpb_inst_2.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAA7FFFF;
defparam sdpb_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAA3FFFFF;
defparam sdpb_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAABFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2AA8FFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAABFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDAAABFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAABFFFFFFFFFFF;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[29:0],sdpb_inst_3_dout[7:6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[13]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 2;
defparam sdpb_inst_3.BIT_WIDTH_1 = 2;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF56FFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF556FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9557FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD556FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5557FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5556FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9555FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD5557FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE5557FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5556FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5555FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFD5557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF5557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF5556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF9555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFD555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFD5557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE5557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFF5556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFF5555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_18 = 256'hFFFFFFFFFFFFEAAAAAAAA5555AAAAA95ABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_19 = 256'hFFFFFFFFFFFE5555555555555555555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1A = 256'hFBFBEFFFFFFFFFFFFFFD5557FFE5555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1B = 256'hBBBFEBFBFFFFFFFFFFF5557FFFD5555557FFEFFFFBBF7EEFBEFFBFFBFBDFEFEF;
defparam sdpb_inst_3.INIT_RAM_1C = 256'hFBBEBFBFFD555555FF5556FFFE5555555FFEFEFFFFF7EFFFFEFBFFFFFEFFFFEF;
defparam sdpb_inst_3.INIT_RAM_1D = 256'hBBFFBFFFFFFE5557F5555FFFF55555557FFFBFFEFF7FBFEFEFFEFFFEFFBBEDFB;
defparam sdpb_inst_3.INIT_RAM_1E = 256'hFBFBFFFFFFF5556FD555BFFF95555555FFFBBFDEF7BBBBFFFFDFEFEFFBEFFFFF;
defparam sdpb_inst_3.INIT_RAM_1F = 256'hBFFFFFFFFFD555FD5557FFFD5555555BFBBEFFEF7BBBBBFBEEFEFFFBFFFFFEEB;
defparam sdpb_inst_3.INIT_RAM_20 = 256'hFFFFFFFFFD555FE5557FFFD55555557FBBEFFFEBFBBFFBBEEFFFFFBFFBFFEFBF;
defparam sdpb_inst_3.INIT_RAM_21 = 256'hFFFFFFFFF555BF5556FFF955555557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_22 = 256'hFFFFFFFF5557F5555FFF955555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_23 = 256'hFFFFFFF9557F9555FFF555555555FFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_24 = 256'hFFFFFFD555FD555BFE555555555FFFFFFAFFFFFFFFFFFFFBFFFFBFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_25 = 256'hFFFFFD555FD5557F9555555555BFFB7EABEDFEEFEBF9BDDFD9F9BF7BEEFFBE9F;
defparam sdpb_inst_3.INIT_RAM_26 = 256'hFFFFE555FF5556955555555557EFDBFF7EDBDEFFEFDFDFBDEFEFFEBFDFFBFDFF;
defparam sdpb_inst_3.INIT_RAM_27 = 256'hFFFF5557F5555AAA555555557EFD7FFBEF7DAFE9FDFDF7E5FFFFEBE9FF7E9FFF;
defparam sdpb_inst_3.INIT_RAM_28 = 256'hFFF5557F5555FFFE55555557EFEBFF7F77EFBFDFDFEF7EFFFFF77FEFF7FEFFFF;
defparam sdpb_inst_3.INIT_RAM_29 = 256'hFF9556FD555BFFF95555557DFBFF67F77EFBD9FDFF6BEFBFBF77E9FA7E9FFFFF;
defparam sdpb_inst_3.INIT_RAM_2A = 256'hFD555FD5557FFFD5555557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2B = 256'hD555FE5557FFFF5555557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h555BF5557FFFF555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2D = 256'h557F5557FFFF555555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2E = 256'h56F9557FFFF555555FFBBBFA7BFDF67DBEBFEDFEAE9E6F77BEBE7A7FFFFFFFF5;
defparam sdpb_inst_3.INIT_RAM_2F = 256'h5FD557FFFF555555FFBFEFFFFFFF7BD7FEFDDFFFFDF7F7BFEBEBFBFFFFFFFF95;
defparam sdpb_inst_3.INIT_RAM_30 = 256'hF955BFFFF555557FFFEEFEBEFFBEBDFE7FEEFFFFAFBFBFEFADFEBFFFFFFFFD55;
defparam sdpb_inst_3.INIT_RAM_31 = 256'hAAAFFFFD55555BFFEDFBFEEFE7EEDADFFEFFFEFFFFFFFEDED9FFFFFFFFFFD555;
defparam sdpb_inst_3.INIT_RAM_32 = 256'hFFFFFF555556FFFDDF7E9DBBEEEEDDDFF6FFDFABEEADADDDEFEFFFFFEAA95556;
defparam sdpb_inst_3.INIT_RAM_33 = 256'h9555555556FFFFFBFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5557F;
defparam sdpb_inst_3.INIT_RAM_34 = 256'hAAAAAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5556AA;
defparam sdpb_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9555AAA;
defparam sdpb_inst_3.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555FFFF;
defparam sdpb_inst_3.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555FFFFF;
defparam sdpb_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF555BFFFFF;
defparam sdpb_inst_3.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5557FFFFFF;
defparam sdpb_inst_3.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9557FFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555FFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555FFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE555BFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5557FFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5557FFFFFFFFFFF;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[23:0],sdpb_inst_4_dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[13],ada[12],ada[11]}),
    .BLKSELB({adb[13],adb[12],adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 8;
defparam sdpb_inst_4.BIT_WIDTH_1 = 8;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'hB1706F6F6F6F6F84FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_04 = 256'h6F6F6F6F6F71FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF56E;
defparam sdpb_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_08 = 256'h6F6F6F6FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7C6E6F;
defparam sdpb_inst_4.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0C = 256'h6F6F70FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD26F6F6F6F;
defparam sdpb_inst_4.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_10 = 256'h6EFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE6E6F6F6F6F6F;
defparam sdpb_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE996F6F6F6F6F6FC8;
defparam sdpb_inst_4.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF76F6F6F6F6F6F76FFFF;
defparam sdpb_inst_4.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF836F6F6F6F6F6FF3FFFFFF;
defparam sdpb_inst_4.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6F6F6F6F6F6FABFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF956F6F6F6F6F72FEFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9716F6F6F6F6FE8FFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD96E6F6F6F6F8FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFEC76D6F6F6F6EFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFEDC6C6E6F6FDAFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFEFBB9D8BACFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3C = 256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_4 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_4_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_9 (
  .O(dout[1]),
  .I0(sdpb_inst_0_dout[1]),
  .I1(sdpb_inst_4_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[2]),
  .I0(sdpb_inst_1_dout[2]),
  .I1(sdpb_inst_4_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_19 (
  .O(dout[3]),
  .I0(sdpb_inst_1_dout[3]),
  .I1(sdpb_inst_4_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_24 (
  .O(dout[4]),
  .I0(sdpb_inst_2_dout[4]),
  .I1(sdpb_inst_4_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(dout[5]),
  .I0(sdpb_inst_2_dout[5]),
  .I1(sdpb_inst_4_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_34 (
  .O(dout[6]),
  .I0(sdpb_inst_3_dout[6]),
  .I1(sdpb_inst_4_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_39 (
  .O(dout[7]),
  .I0(sdpb_inst_3_dout[7]),
  .I1(sdpb_inst_4_dout[7]),
  .S0(dff_q_0)
);
endmodule //Gowin_SDPB2
