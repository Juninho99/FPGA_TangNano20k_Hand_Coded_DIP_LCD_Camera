//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Sat Aug 12 15:43:55 2023

module Gowin_SDPB1 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);//sobel_3x3

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [14:0] ada;
input [7:0] din;
input [14:0] adb;

wire lut_f_0;
wire lut_f_1;
wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [1:1] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [2:2] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [3:3] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [4:4] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [5:5] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [6:6] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [7:7] sdpb_inst_7_dout;
wire [29:0] sdpb_inst_8_dout_w;
wire [1:0] sdpb_inst_8_dout;
wire [29:0] sdpb_inst_9_dout_w;
wire [3:2] sdpb_inst_9_dout;
wire [29:0] sdpb_inst_10_dout_w;
wire [5:4] sdpb_inst_10_dout;
wire [29:0] sdpb_inst_11_dout_w;
wire [7:6] sdpb_inst_11_dout;
wire [27:0] sdpb_inst_12_dout_w;
wire [3:0] sdpb_inst_12_dout;
wire [27:0] sdpb_inst_13_dout_w;
wire [7:4] sdpb_inst_13_dout;
wire [23:0] sdpb_inst_14_dout_w;
wire [7:0] sdpb_inst_14_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire mux_o_6;
wire mux_o_8;
wire mux_o_16;
wire mux_o_18;
wire mux_o_26;
wire mux_o_28;
wire mux_o_36;
wire mux_o_38;
wire mux_o_46;
wire mux_o_48;
wire mux_o_56;
wire mux_o_58;
wire mux_o_66;
wire mux_o_68;
wire mux_o_76;
wire mux_o_78;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_0.INIT = 16'h4000;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_1.INIT = 16'h4000;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8B6FFFFFFFFFFFFFFFFE;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7B3FFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFFFFFFBF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB5;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFDFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFF3FC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FEBFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFF5FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFC9FFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFF7FF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFDFFF;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFF7FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFDFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFDFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA7FE7FFFFFF;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hFFFFFFE7FF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3F;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFDFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF7FFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF9FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FE3FFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFC7F;
defparam sdpb_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFF3FF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFEFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hFFB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFDFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFEBFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFE7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF9FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFE3FFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_22 = 256'hFFFE7FF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF0F;
defparam sdpb_inst_0.INIT_RAM_23 = 256'hFFFFF7FFFFFFEFFD7FFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFF3FFFFFFB59FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFE00000003FFF00027F8BFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_26 = 256'hF77FFF1FABFFFFF7BFBFEFADA9066FD8000000FFFC0027FF02BFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_27 = 256'hFFE4FFEB5B73FFEEDF5F3F66DD87CBBBE23D5BFA0000003FFF804FFFFEA9FF8C;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h7FF7FFD7FFFF13F856A3BFF0B7ABFBB054B3848AFCE898FD7FFFFFFBFFD00DFF;
defparam sdpb_inst_0.INIT_RAM_29 = 256'hFFFFFFFFCFFFFFF3FFFFFFFEBBFE1F34BEE7FF3EFAFEDDFFF3B7B33FFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2A = 256'hF81D53B7FE000003FFFFDFF5FFFFF4FFBB3FFBC1175F9FC7BF67FBA8E1F47E8F;
defparam sdpb_inst_0.INIT_RAM_2B = 256'hFD664BCFF0592DDEBFEFF7FEAFBFE3FF8FFFFFEFE747F977FDC4FF71EFCFFEF6;
defparam sdpb_inst_0.INIT_RAM_2C = 256'hF19C28F1BE6BAE63544E6F53EFF800E7D31FFFFFFBFFFFFFFAD9F19C3BB0ABEB;
defparam sdpb_inst_0.INIT_RAM_2D = 256'hFFEBCDF3C31D05BC9FDFDFC8EAFF98BFA7FA00FE1AF3FF3FFEFFFFFF7FFFFCAF;
defparam sdpb_inst_0.INIT_RAM_2E = 256'hFFC7FFFFF3FB57F6F1E54DB74FEBE377DF9A665FD1FFFFF7FF7DFFF3FF7FFFFF;
defparam sdpb_inst_0.INIT_RAM_2F = 256'hDFFFEFFEFFF9FFFFFE7E9B7F067D92AFE67FFADEF1A3B9BEBEFFFFF5FFFFBFFE;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h3B57FFFFF7FEADFFDFFF7FFFFFE7F0BF2492CCBE3E7EBB7ED887824E6E7FFFFF;
defparam sdpb_inst_0.INIT_RAM_31 = 256'hCDFF7FF7F31CFFFFFCFFFFBFF7FFDFFFFFF7E8E7048729BA3FDFECCAD83EC748;
defparam sdpb_inst_0.INIT_RAM_32 = 256'hA0F2FEFF973DB1D5EBECFFFFFCFFE75FFF7FFFFFFFFFFFEB3DFF6BAF3FFDFFFF;
defparam sdpb_inst_0.INIT_RAM_33 = 256'hFF17FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FCF7FFEFFDFFFFFFBFF68F2967D6;
defparam sdpb_inst_0.INIT_RAM_34 = 256'hFFFFFB7FFFEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFEFFFFFEFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_35 = 256'hEFFFFFC7FFFFFEDF9BBBFF9FF7FFDF7FDFFFFDEBFFF7FEFFFFFEFFCE3FFDFFBF;
defparam sdpb_inst_0.INIT_RAM_36 = 256'hFFFFFFFC65FFDFEFFFFFFFDD751D73A3D9E7B71B1FAB3D47DF7C77BFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h3F1FD797FFFFFAFF3B7FF6DCFFFFFFFBF847C794FF1C5C7FC1D56942FC8E9D6F;
defparam sdpb_inst_0.INIT_RAM_38 = 256'hFF1A9FBEAB7BF9FCFFFFFEDFF9DFFFBCFFFFFFFFF359E262FF879BD5E2E4DE7D;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h9EF8777D7D0FFBFFECECFE7F7FFFFFEFFDFFFFDEBFFFFFFFBBF9F91CCF7DFBFD;
defparam sdpb_inst_0.INIT_RAM_3A = 256'hF9BFE7AED8337C4F9FB0E5FFEEB0CFFE5FFFFFEBFFFD7FFE3FFFFFFFFFFEBD46;
defparam sdpb_inst_0.INIT_RAM_3B = 256'hA7E7FFFFFFF7A8D77B3FFF03F7DD323EFF9C1FFF83FFFFFF7FEF9FFDC07FFFFF;
defparam sdpb_inst_0.INIT_RAM_3C = 256'hFBFF4FFFEFFF5FFFFF9D67FCCF27B9FCF9EB6E6FCFA7FDF87E7FFFFFFFFFEFFF;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h8EF7FFFFFEFFC77FFBFFB3FFFFF76B6DB7D9D6F87E7E670FF7B4C071304FFFFF;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h5FB934EFE9B4FFFFFFBFFFD7FE7FD1FFFFFDC3BB30FA8E9C5FAFC9E4FBFF1B39;
defparam sdpb_inst_0.INIT_RAM_3F = 256'hFFFFFDCDF7FFE7FEDFFFFFFFFFFFFEFFFFD7FF5FFFFFF6DFF4FA3F7B9FE7FE76;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F7FFFFFFFFFFFFFFFFE;
defparam sdpb_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE3FFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_02 = 256'hFFFFFF7FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFEFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFBFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FCFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3FFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_08 = 256'hFFBFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFBFF;
defparam sdpb_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFEFFEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0F = 256'hFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFBFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFBFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_15 = 256'hFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFF;
defparam sdpb_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFDFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFF3FFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFDFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1B = 256'hFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hFFFFFFFDFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3;
defparam sdpb_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF7FF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFEFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_22 = 256'hFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF7F;
defparam sdpb_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFD1DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFF00000001FFF0001FFE1FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_27 = 256'hFFF8FFFEDFFDFDEFEF9F7F6ED9D1FAF7CBA26FE80000002FFFFF9FFFFF1FFFFF;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h7FFFFF7FFFFF5FFDD77FBD71FBEFCCE96C8F7CBA594D9DFE7FFFFFFDFFFFF5FF;
defparam sdpb_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFEFFFFFDBFF79DEDFDCFDF5FB7EFEDFDE7726F3D7BFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2A = 256'hF96F9D6FFEFFFFFFFBFFDFFDFFFFFF7F9B779BE3271BBFDFDF33F79BD7B2E74F;
defparam sdpb_inst_1.INIT_RAM_2B = 256'hFBC7F9BD78597E5FFF9FFF9FBEFFFFFF9FFFFFCFFFEDFAFACEC7EFFBE7FFFC57;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h56B4BBF7BE72EFEB2E7B698BBFF7FDFFE7CFFFFFFFFFFFF9FFFBE29ED3B055EF;
defparam sdpb_inst_1.INIT_RAM_2D = 256'hFFFED7EFE7FFA5FF7FFFBDFEC877DF956FFDFFFFFFF7FF7FFFFFFFFF7F757CBF;
defparam sdpb_inst_1.INIT_RAM_2E = 256'hFFF7FFFFF7FBF7F25687D3BFDDFBE7F3FF3CF6DCB9FFFFFFFF7DFFFFFFBFFFFF;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h7FFFCFFFFFFBFFFFFF7ECFFFF1FB9A4DFFFEF9FDF0FFB5DFBEFFFFFFFFDF7FFB;
defparam sdpb_inst_1.INIT_RAM_30 = 256'hFAAFFFFFE7FEFFFFFFFEFFFFFFDF81DD18F976E97F1FB8B3743ADF6D7D1FFFFF;
defparam sdpb_inst_1.INIT_RAM_31 = 256'hF7FFFFFFFFFFFFFFFDFFB8BFFFFFBFFFFFFBF17F4E67DF7BDFEFFE9CCC37E3DC;
defparam sdpb_inst_1.INIT_RAM_32 = 256'hFFFF7F7FEFF7FFBFFFFFFFFFFF7FFF9FFDFFEFFFFFFF7FFEFEFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_33 = 256'hFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFEFFF9FFFFFFFFFBFEFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFD1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFE7FDFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hFFFFFFF7FFFFFF7EFFFF7F7FFFFFFFFFFFFFFFFF7FFDBFFFFFFF7FFBFFFFFF3F;
defparam sdpb_inst_1.INIT_RAM_36 = 256'hFFFFFFFF7FFFDFE7FFFFFFFE655F3FDFFFFFF7FE3FBB7FAFEF7C7FBFFFFFDFFA;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h5FDF9FE3FFFFFDFFAF7FFBBFFFFFFFF98EDFF3D4773C2EFF77D3DD2A7C3F9E0F;
defparam sdpb_inst_1.INIT_RAM_38 = 256'hE7DDC7DFAFF1FDFCFFFFFFFFF3DFFFFFFFFFFFFF77E7E5F98CC76FFDD3E1B51F;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h89F1F9FC78FFA7FFFDD07FF8FFFFFFFFFFFFFF9FFFFFFFFFFCF5F9BF937DF9FB;
defparam sdpb_inst_1.INIT_RAM_3A = 256'hFFBF9FFBE97ADC3FFF1FE2FDFC3E5FFF4FFFFFFFFFDCFFFA37FFFFFFEEBF7D73;
defparam sdpb_inst_1.INIT_RAM_3B = 256'hE7EFFFFFFFF7D5FFF81E9743F78F7DBEFC8F1FE1CBFFFFFF7FEFBFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3C = 256'hF7FF7EFFF003FFFFFFDFFDB39FAFBDFDFFFBFEFFFF97FFF8FF7FFFFFDFFFE7FF;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h3703FFFFFEFFCF3FFBFF87FFFFF7FFDF7BEFFF7FBF7DCF77E7FF7EFE3FDFFFFF;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h1FBFEFD3ABFDFFFFFFBFF9F7FF7FFBFFFFFDEEBF86F679BCBFEF95CEFDED18EC;
defparam sdpb_inst_1.INIT_RAM_3F = 256'hFFFFFDFFBFFFFFFFFFFFFFFFFFDFFE6BFFFFFF1FFFFFF3CEF7FBBFF35FE3F3F9;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE6C7FFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_02 = 256'hFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_2.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFCFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFBFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FD3FFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFF;
defparam sdpb_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFBFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF9FFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFF;
defparam sdpb_inst_2.INIT_RAM_0F = 256'hFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFDFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF7FF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_15 = 256'hFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF;
defparam sdpb_inst_2.INIT_RAM_16 = 256'hFFFFFFFFFFFDFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1B = 256'hFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1C = 256'hFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF5F;
defparam sdpb_inst_2.INIT_RAM_23 = 256'hFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFF7FFFFFFF53FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFD0079FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_27 = 256'hFFFFFFFFBD7DFFFBDFFFFF70F9D9F7F2EF3677FDFFFFFFDFFFFFFFFFFF8FFFFF;
defparam sdpb_inst_2.INIT_RAM_28 = 256'h7FFBFF7FFFFFDFFFD7C33DFDF7D7EFEA058E9BB67CDE19FE7FFFFFFBFFEFFFFF;
defparam sdpb_inst_2.INIT_RAM_29 = 256'hFFFFFFFFDFFEFFEFFFFFD7FF63FF6F7CBD677BFE7FDDDE77A7BFF77FFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2A = 256'hFD3FFB33FFFFFFFFF3FF9FFFFFFFFFFFB97FB7DBBF5D9ECFFFB3B39BFBF6FCCF;
defparam sdpb_inst_2.INIT_RAM_2B = 256'hFFE3DBFF58F976EFFFBFFF9F7CFFF7FFFFFFFFFFF7FFF870ECC7E73BEFCCFDEF;
defparam sdpb_inst_2.INIT_RAM_2C = 256'h668CFEFFBEFAEEF7345B6BDFBFF7FFFFF7AFFEFFF7FFFFFFFFDBE59D1971FFCE;
defparam sdpb_inst_2.INIT_RAM_2D = 256'hCFDCEFC9D3BB96FE67BFFBBFDDFF5B53EFFE00FFFDE7FFBFFFFFFFFF7FFBFC77;
defparam sdpb_inst_2.INIT_RAM_2E = 256'hFFE7FFFFF3FBFDF7F02FC1B7DFFFE7FFB3FFE6779DFFFFE7FF7DFFEFFF3FFFFF;
defparam sdpb_inst_2.INIT_RAM_2F = 256'hFFFBFFFFFFFBFFFFFF7EF47DB879F3EFFF7DFFDFFEFF71F3377FFFFDFFEF7FFD;
defparam sdpb_inst_2.INIT_RAM_30 = 256'hFF67FFFFFFFEFFFFDFFFFFFFFFFFC79D1B9FECE23C9F7133F4FFEC656CFFFFFF;
defparam sdpb_inst_2.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFEBFF7FFFFFFFFFFF3F7B78E59BF6F6FED2EF8EF8FDB;
defparam sdpb_inst_2.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFDFFFFFEFFFFFFF7FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_33 = 256'hFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF7FFBFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFBFFFE7FEFFFFFFF7FF;
defparam sdpb_inst_2.INIT_RAM_35 = 256'hFFFF7FD7FFFFFFBFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFF3F;
defparam sdpb_inst_2.INIT_RAM_36 = 256'hFFFFF7FFFFFFFFF7FFFFFFEEF7DE9F37FCFF77BFBF3F7FF9EFFEF7BFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_37 = 256'hDEE7F7FBFFFFFDFFBFFFFFFFFFFFFFFB8FB74BC4FFDE3E1F87C2D17A7C5F1E0F;
defparam sdpb_inst_2.INIT_RAM_38 = 256'hE73F9FFFD3F3FBFDFFFFFFFFFBFFFEFDFFFFFFFF7FBFDFF6FEFFE79FF5FC3B7E;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h59CA79FF7DC72FE7F2E17E78BFFFFFEFFEFFFFDEFFFFFFFFDCFD71FCBF7DFAF7;
defparam sdpb_inst_2.INIT_RAM_3A = 256'hFDAFBFFEFBF85C2F9F77D1FDFFBA3FDE2FFFFFFFFFBCFFFAF7FFFFFFEE7E9FE7;
defparam sdpb_inst_2.INIT_RAM_3B = 256'hD81FFFFFFFF3FDFFB8FFFFE3F7BE7CFF7F2FEFEFF3FFFFFEFFFFBFFE3FFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3C = 256'hFFFFFFFFE005FFFFFFDCFC3BDE2799FFFBE3BD5FCF8FF9FEFDFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3D = 256'hBEFFFFFFFEFFEFBFFBFFD7FFFFF77EEE7FA9EEFFFEFEFF77EFF7FF7F7F9FFFFF;
defparam sdpb_inst_2.INIT_RAM_3E = 256'h1F3EE7B3D7C9FFFFFFFFFBE7FF7FFFFFFFFDEF3BADEFFDDCDFCF8BE7FFF97FAD;
defparam sdpb_inst_2.INIT_RAM_3F = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFF7FFFFFFDFFFDFFFFFF1CFF8789EABA3F3F9F5;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8DBFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_3.INIT_RAM_01 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEF7FFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_02 = 256'hFFFFFF7FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFEFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FD7FFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_08 = 256'hFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF;
defparam sdpb_inst_3.INIT_RAM_09 = 256'hFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFBFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0F = 256'hFFFFFFF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF;
defparam sdpb_inst_3.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFEFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF;
defparam sdpb_inst_3.INIT_RAM_16 = 256'hFFFFFFFFFFFDFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFF7FFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFBFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1B = 256'hFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1C = 256'hFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE7FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF9FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_22 = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5F;
defparam sdpb_inst_3.INIT_RAM_23 = 256'hFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFF7FFBFFFE6BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFDFFF5FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_27 = 256'hFFF9FFFFBD8DFBF5DFDFFF9B364E3CCCF5FF77FBFFFFFFFFFFFFFFFFFFAFFFFF;
defparam sdpb_inst_3.INIT_RAM_28 = 256'hFFFBFF7FFFFFDFFFEF41FFFBF78FDCD60FE11C63FCFC9DFE80000007FFFFFBFF;
defparam sdpb_inst_3.INIT_RAM_29 = 256'hFFFFFFFFDFFEFFE7FFFFDBFFFDFFFFBDDEFFFB3FFFDE9E7FA75FD33FFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_2A = 256'hFD76DBF3FFFFFFFFF3FFDFFCFFFFFFFFB93FD3E7FF9BDECFDF77F7DFE7D6CDEF;
defparam sdpb_inst_3.INIT_RAM_2B = 256'hFDFB9F9F57C9AEFEFFBFFF9F3EFFF7FFBFFFFFDFEF6FFFF9DCFFFF3BF7CCEDE7;
defparam sdpb_inst_3.INIT_RAM_2C = 256'hB6FF37FDBEF7E7FF4FDB6D73FFFFFFFFE7EFFDFFFFFFFFFDFBFBEFDE9CFFFDCF;
defparam sdpb_inst_3.INIT_RAM_2D = 256'hFFEEEFDFE2FF86FE67CF9BBCEDF75FF27FFFFF3FFDF7FF3FFDFFFFFF7F7F7B6F;
defparam sdpb_inst_3.INIT_RAM_2E = 256'hFFE7FFFFF3FB35F6FA67D1B7BFFBF77BDF3DC7F4FFFFFFFFFF7DFFFFFF7FFFFF;
defparam sdpb_inst_3.INIT_RAM_2F = 256'hFFFBFFFF7FFBFFFFFFFFFF7F5EFBB71CF77FF9DEF7EF75F9AF7FFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_30 = 256'h5B0FFFFFFFFFFFFFFFFFFFFFFFDFDF9EBF3FF5DFFFBFFEF3EE734D7DFEDFFFFF;
defparam sdpb_inst_3.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFDFFDEBFF7FFFFFFFFFBFFFF766EFBFA0FDFECEEDBCFFBBF;
defparam sdpb_inst_3.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7FF7FFFEFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_33 = 256'hFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEF7FFFFFBFFFFFFDFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_34 = 256'hFFFFFDFFFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFBFFFF7FEFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_35 = 256'hEFFF7FD7FFFFFFBFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFF7F;
defparam sdpb_inst_3.INIT_RAM_36 = 256'hFFFFFFFF7FFFFFF7FFFFFFFEF9BF7F73FDF0F07F3FC783DBF0FFF07FFFFFDFFD;
defparam sdpb_inst_3.INIT_RAM_37 = 256'h5F2FF78FFFFFFDFFBEFFFFFBFFFFFFF99E0FBFFD73FFFFEF77DDCE6FFF9F7DFF;
defparam sdpb_inst_3.INIT_RAM_38 = 256'hF37FBFBF9FF9FFFDFFFFFF7FF7FFFEFFFFFFFFFF7BFFE4F5DDD70B3386FB31BD;
defparam sdpb_inst_3.INIT_RAM_39 = 256'h75D6F1FFF9CFBBF7E2F3FE787FFFFFEFFFF7FFFFFFFFFFFFFCF6F55CB7F1FBFF;
defparam sdpb_inst_3.INIT_RAM_3A = 256'hFDFFF7FAF0FBDDEFDE7FD1F9FDF9FF9FFFFFFFFBFFFEFFF3F7FFFFFFEEFFBFE7;
defparam sdpb_inst_3.INIT_RAM_3B = 256'hFFFFFFFFFFF3F7FEFADF1F43FF9D7BBEFEBF07FF8FFFFFFE7FFFBFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3C = 256'hFFFF7FFFF003FFFFFFDFF0B98E7FFBFCFBFB7FEFBFD3FDFEFFFFFFFFFFFDFFFF;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h2F1FFFFFFFFFEFBFFBFFD7FFFFF77D6FEFBFE6FFBE7F7753EFEFFEFE3FDFFFFF;
defparam sdpb_inst_3.INIT_RAM_3E = 256'h7EFEDFFBFBFFFFFFFFFFFFD7FF7FFFFFFFFDCFFFB5FAFDDE0FDFA3CFFEF7DA3E;
defparam sdpb_inst_3.INIT_RAM_3F = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFF7BFFFFFFDFFFFFFDFCF67FFE6FFFF3FFF5;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF937FFFFFFFFFFFFFFFFE;
defparam sdpb_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF117FFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_02 = 256'hFFFFFF001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01;
defparam sdpb_inst_4.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFE007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC02FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF802FFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_08 = 256'hFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFF;
defparam sdpb_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFE000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0E = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0007FFFFFF;
defparam sdpb_inst_4.INIT_RAM_0F = 256'hFFFFFFE8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam sdpb_inst_4.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFE002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0013FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_15 = 256'hFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001FF;
defparam sdpb_inst_4.INIT_RAM_16 = 256'hFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC002FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4003FFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1B = 256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFF;
defparam sdpb_inst_4.INIT_RAM_1C = 256'hFFFFFFFE000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam sdpb_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_22 = 256'hFFFE0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00BF;
defparam sdpb_inst_4.INIT_RAM_23 = 256'hFFFFFFFFFFFF9000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFF8007FFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFF7FFFFFFE000FFFE003FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000001FFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_27 = 256'h0005FFEEFF0FFBF3FFBF778610787987FFFBFFF80000000000000000005FFFFF;
defparam sdpb_inst_4.INIT_RAM_28 = 256'h0003FF4000003FFFDF617E7CFB83DDDE8DFF1E21B97EDFFFFFFFFFF800100800;
defparam sdpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFC001FFF800002BFFE7DEEFDCDDECF7FEFCFE9E7F6E5BF7FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2A = 256'hFDA699F3FFFFFFFFF4003FFF000000FFFFF797FBB77B9CDFBFB3B799EB9BC6FF;
defparam sdpb_inst_4.INIT_RAM_2B = 256'hFDC7FFFF187D3DDFFFC000603F000FFF8000002FE76DFFFFCCDFEF3BE7CFECEE;
defparam sdpb_inst_4.INIT_RAM_2C = 256'hE79DFFFFFF79FF77CE3A6FFFBFF000001FD001FFF0000007FDDF60FFB8F6FBFE;
defparam sdpb_inst_4.INIT_RAM_2D = 256'h0FFCD7D9FDDFEEFE67FFFBFEFDF61BF2FFFFFF0001F800FFFE0000007FB358EF;
defparam sdpb_inst_4.INIT_RAM_2E = 256'hFFE800000BF333FB7EF6D5BFFDFBEF7FBBBFD7E6BBFFFFE0007E001FFFC00000;
defparam sdpb_inst_4.INIT_RAM_2F = 256'h8003C000FFFC0000007EFFFFDBED974DF6FDFBDEECCF7D97E7FFFFFE001F8003;
defparam sdpb_inst_4.INIT_RAM_30 = 256'hFB9FFFFFF000F8001FFE0000002F9F9C73FFFDFBBCFFB877A2FA1F646EFFFFFF;
defparam sdpb_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFE001F4007FF80000003F9F77E2F7DFB3F87EFFCEBEFBFFF;
defparam sdpb_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF800FA001FFE0000000FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_33 = 256'hFF97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001F0003FF80000001FFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_34 = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007C001FFE0000000FFF;
defparam sdpb_inst_4.INIT_RAM_35 = 256'hE000FFE80000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FC003FFC0;
defparam sdpb_inst_4.INIT_RAM_36 = 256'hFFFFF80078000FF00000000F7BBF9FBBCEF0783F3F87839DE0FEF87FFFFFC003;
defparam sdpb_inst_4.INIT_RAM_37 = 256'h7ED7EFF3FFFFFC005F0007FC00000007DFE7C3FCFF7C1E1F0FC0C0E6F87F9E1F;
defparam sdpb_inst_4.INIT_RAM_38 = 256'hEB7DEFFFA7F5FBFFFFFFFF800FC001FE000000006F8BD9FF1CDF674FE9F3BE5C;
defparam sdpb_inst_4.INIT_RAM_39 = 256'h9DE3787E7BF77FEFF2F2FE783FFFFFE000F0003E000000001FF071FD0FBFF8F3;
defparam sdpb_inst_4.INIT_RAM_3A = 256'h03DF87F9E87C1C1FFEF3EEF9FC3C1FDF1FFFFFFC007E000408000000173FBEFF;
defparam sdpb_inst_4.INIT_RAM_3B = 256'h0000000000F3E3FF389F07CBEFEEF43FFE0F0FE7C3FFFFFF800F800000000000;
defparam sdpb_inst_4.INIT_RAM_3C = 256'hF0007C0010040000001EFF7BEEFFBFFFF9FF9EDF9FE3F9FDFCFFFFFFE003E000;
defparam sdpb_inst_4.INIT_RAM_3D = 256'h1F0FFFFFFE000FC007FFA8000007BC4F73DDF6FF3FFFEF13F3EEFE7EBFBFFFFF;
defparam sdpb_inst_4.INIT_RAM_3E = 256'hBE7FE7078381FFFFFF8007C800FFFC000001DFBBC3E7FFDD3FFFB5DEFCF13E1E;
defparam sdpb_inst_4.INIT_RAM_3F = 256'hFFFFFE7FFFFFFFFFFFFFFFFFFFF001F8003FFFA00000FBCDF97D9E7707EFF1F3;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b0;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDE7FFFFFFFFFFFFFFFFE;
defparam sdpb_inst_5.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_02 = 256'hFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE;
defparam sdpb_inst_5.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFBFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEFFF;
defparam sdpb_inst_5.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0F = 256'hFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF;
defparam sdpb_inst_5.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_15 = 256'hFFF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFBFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;
defparam sdpb_inst_5.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_22 = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFF;
defparam sdpb_inst_5.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_27 = 256'hFFFDFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_28 = 256'h7FFBFFFFFFFFBFFBE7FBFF77F387DDE4FE97EBADB9FCDDFF00000003FFEFF7FF;
defparam sdpb_inst_5.INIT_RAM_29 = 256'hFFFFFFFFDFFEFFFFFFFFFFFFE5FEEFFFFFFFFFBEFDCF9FFFEE5FF77FFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2A = 256'h7B66F53FFFFFFFFFFFFFFFFFFFFFFF7F9FBFDBFFF79FFDFFFFBFFFFFFD96EFEF;
defparam sdpb_inst_5.INIT_RAM_2B = 256'hF9C3FDDF9979EF7EFFFFFFFF7FFFFFFFBFFFFFFFFFFFFFFEEFFFF7BFEFFFFEF6;
defparam sdpb_inst_5.INIT_RAM_2C = 256'hF7EFBDFFFF70F6F7F63E7DFBFFF7FFFFFFFFFDFFF7FFFFFFFFFFF1BFBDFFFFEF;
defparam sdpb_inst_5.INIT_RAM_2D = 256'hEFECDFFDFFDB6EFFEFFFFFFDCDFE1F7EFFFFFFBFFDFFFFFFFDFFFFFFFFFEFCA7;
defparam sdpb_inst_5.INIT_RAM_2E = 256'hFFEFFFFFFBFBBBFBED67E9FBBBF7E7FFF37DC7F4D9FFFFFFFF7DFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2F = 256'hBFFFFFFF7FFFFFFFFFFFFEFFDFFFBF6EFFFDFDFFFFCFB595FEFFFFFDFFEFFFFF;
defparam sdpb_inst_5.INIT_RAM_30 = 256'hBBCFFFFFEFFEFBFFFFFEFFFFFFFFD79F9AFD6FD9FEBFFFFF3EFFDF77FDFFFFFF;
defparam sdpb_inst_5.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFDFFFEFFF7FFBFFFFFFBF8FF873FFFFB9FCFEE1DEC7F87DD;
defparam sdpb_inst_5.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7FF7FFFEFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_33 = 256'hFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFBFFFFFFFFFDFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_34 = 256'hFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBDFFFFFEFFFFFFF7FF;
defparam sdpb_inst_5.INIT_RAM_35 = 256'hFFFF7FDFFFFFFFBFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFF;
defparam sdpb_inst_5.INIT_RAM_36 = 256'hFFFFF7FF7BFFFFF7FFFFFFEFFFFF3FFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFDFFF;
defparam sdpb_inst_5.INIT_RAM_37 = 256'hBEFFF77BFFFFFDFFDFFFFFFFFFFFFFFFDEF7BBFFF3FFFFFF7FFFFFFEFBFFFFEF;
defparam sdpb_inst_5.INIT_RAM_38 = 256'hFBFEEFDFFFFFFBFFFFFFFFFFFFFFFEFDFFFFFFFFEFFFF1F7FCDF7FFFE6FBFFFD;
defparam sdpb_inst_5.INIT_RAM_39 = 256'hFDF3FEBFFEDF7FEFF7FD7FFF7FFFFFFFFEFFFFFEFFFFFFFFDBFCFFFFF777FFFF;
defparam sdpb_inst_5.INIT_RAM_3A = 256'hFDEFB7FBF6FFFFEFDFBDD3FFFDBFDFDFEFFFFFFBFFFEFFF87FFFFFFFFFFFDFFF;
defparam sdpb_inst_5.INIT_RAM_3B = 256'hFFFFFFFFFFF3E7FEF83F97CBEFEF7FFFFFFF0FEF8BFFFFFFFFF7FFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3C = 256'hFFFF7DFFEFFBFFFFFFDDFFF9BF67BBFFFDFFDD6FBFFBFFFBFFFFFFFFDFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3D = 256'h2E17FFFFFEFFFFFFFFFFDFFFFFF7BDFE7FEDEF7F7FFFD7F3EFEFFE7FFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3E = 256'hFFBDDFFF7BFDFFFFFFFFFBFFFF7FFBFFFFFDDFBBEFEEF9DF2FFFB7F5FBFD7E3C;
defparam sdpb_inst_5.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFBFFDFFF7FFFFFF7ADF7FAFF6FFFEFEFFD;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[6]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b0;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDEFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_6.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_02 = 256'hFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE;
defparam sdpb_inst_6.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFBFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_09 = 256'hFFFFFFFFFFEFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFF;
defparam sdpb_inst_6.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_15 = 256'hFFF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF;
defparam sdpb_inst_6.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1C = 256'hFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFBFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDF;
defparam sdpb_inst_6.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFF7FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFDFFFFF;
defparam sdpb_inst_6.INIT_RAM_28 = 256'h7FFFFFFFFFFFBFFBFF437FFC77D7DDE58C9B1E30BF6EDDFFFFFFFFFFFFFFFBFF;
defparam sdpb_inst_6.INIT_RAM_29 = 256'hFFFFFFFFFFFEFFFFFFFFFFFEFDDF5FDDDDEFF77EFDFEFEFFFFDB777FFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2A = 256'hFB7DB7FBFFFFFFFFFFFFFFFFFFFFFFFFFD77DBF7777FBFEFBF7BB7BBFDF6DDDF;
defparam sdpb_inst_6.INIT_RAM_2B = 256'hFFFBFBBCFEEFB56EFFBFFFFF7FFFF7FFFFFFFFFFF76DFFFEFDD7EFFBFFEFEEF7;
defparam sdpb_inst_6.INIT_RAM_2C = 256'hFF8DBDFFBF7EEF77C7DBED7BBFF7FFFFFFBFFDFFF7FFFFFFFFDB7DBFFB35F7EE;
defparam sdpb_inst_6.INIT_RAM_2D = 256'hFFDFD7EFF3BB0DFEFFFFBDFEFDF7FB56EFFFFFBFFFFFFFFFFFFFFFFF7FF75F7F;
defparam sdpb_inst_6.INIT_RAM_2E = 256'hFFEFFFFFFBFFBDFB7FBEDF7FDDF7FF7FBF7DDEDFBFFFFFFFFF7DFFEFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2F = 256'hBFFBFFFFFFFBFFFFFF7EFE7FDBEDF77EF7FEFDDDFEFF7BFBB77FFFFFFFFF7FFF;
defparam sdpb_inst_6.INIT_RAM_30 = 256'hBF8FFFFFFFFEFBFFDFFFFFFFFFFFBFDFB6FB75EB3DFFBFF7FDFBEFF7ED9FFFFF;
defparam sdpb_inst_6.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFDFFFFFFF7FFFFFFFFFFF1F70E6F5D7F1F8FFE1FF82EC3BD;
defparam sdpb_inst_6.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFBFFBFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_34 = 256'hFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFEFFFFFFF7FF;
defparam sdpb_inst_6.INIT_RAM_35 = 256'hEFFF7FFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_36 = 256'hFFFFF7FFFFFFFFF7FFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFF;
defparam sdpb_inst_6.INIT_RAM_37 = 256'hFF1FFF8FFFFFFFFFDFFFFBFBFFFFFFFF9EFFBFDDF37FFDFFF7DFFFFBFBFFFDFF;
defparam sdpb_inst_6.INIT_RAM_38 = 256'hFF7FFFFFBFFFF9FEFFFFFFFFFFDFFEFFFFFFFFFFFFEDF5FFFEFF8F93EBF8F93F;
defparam sdpb_inst_6.INIT_RAM_39 = 256'hEFFDFFFFFFFF3BE7F3FFFE7F3FFFFFEFFFFFFFFFFFFFFFFFFFFE7FDFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3A = 256'hFDFFF7FFF87FFFFFFFFFF2F9FDFFFF9FEFFFFFFFFFFEFFF77FFFFFFFF7FE9FEF;
defparam sdpb_inst_6.INIT_RAM_3B = 256'hFFFFFFFFFFF7E7FFFA9F7FBFE7FFFFBEFFAFE7FFF3FFFFFFFFFFBFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3C = 256'hFFFF7DFFEFFDFFFFFFDCFDFFFE6799FEF9FBFFCFFFB3F9FFFFFFFFFFDFFDFFFF;
defparam sdpb_inst_6.INIT_RAM_3D = 256'h3E1FFFFFFEFFFF7FFFFFDFFFFFF73FFE6FA9E67F3EFDFFFBFFEDFF7FFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3E = 256'hFFFDFFFFFFBFFFFFFFBFFBFFFFFFFBFFFFFDFFBFE7FBF99F2FBFA7FFFFFFFE3E;
defparam sdpb_inst_6.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFFF7FFFFFFFFCFFFFFE7FFFFFFEFF;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[7]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b0;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1FFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_02 = 256'hFFFFFF803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE01;
defparam sdpb_inst_7.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFF003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_08 = 256'hFF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFF;
defparam sdpb_inst_7.INIT_RAM_09 = 256'hFFFFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0E = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0F = 256'hFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sdpb_inst_7.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_15 = 256'hFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001FF;
defparam sdpb_inst_7.INIT_RAM_16 = 256'hFFFFFFFFFFFE000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1B = 256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFFFFF;
defparam sdpb_inst_7.INIT_RAM_1C = 256'hFFFFFFFE000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam sdpb_inst_7.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFC003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_22 = 256'hFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003F;
defparam sdpb_inst_7.INIT_RAM_23 = 256'hFFFFFFFFFFFFC001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFF800000000000000001FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000007FFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_27 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000003FFFFF;
defparam sdpb_inst_7.INIT_RAM_28 = 256'h8007FF8000007FFFBFFFFEFBFFFFFFFBF77EFDFFFFFFFFFFFFFFFFFC001FFC00;
defparam sdpb_inst_7.INIT_RAM_29 = 256'hFFFFFFFFE001FFF0000007FFFFFFFFBFFEFEFFFFFFFFFFEFBFFFBFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFF8003FFE000000FFFFFFFFEFFFFFFFFFFFFFFFFFEFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2B = 256'hFFFFBFFFFFFFFFFFFFC00000FE000FFFC000001FFFFFF6FBFFFFFFFFFFFEFFFF;
defparam sdpb_inst_7.INIT_RAM_2C = 256'hBF7FFBFBFFFFFFFFBFFFFFDFFFF800000FC003FFF8000003FDFFFFFEFFFFFBFF;
defparam sdpb_inst_7.INIT_RAM_2D = 256'h1FFFFFFFEDFFFFFFFFDFFFDFFFFFFFFFFFFFFFC003F0007FFE000000FF7FFFFF;
defparam sdpb_inst_7.INIT_RAM_2E = 256'hFFF0000007FFFFFFFBFFFFFFFFFFFFF7FFFFFFFFFFFFFFF000FE001FFF800000;
defparam sdpb_inst_7.INIT_RAM_2F = 256'hC007E000FFFC000000FFEFFEFEFFFFFFFF7FFFFFF7FFFFFFFFFFFFFE001F8003;
defparam sdpb_inst_7.INIT_RAM_30 = 256'hFFFFFFFFF001FC003FFF0000001FFBFFFFBFFFFFFFDFFF7FFFBFFEFEFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFE003F000FFFC0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF800FC001FFF0000000FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE001F8007FFC0000003FFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_34 = 256'h000001FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC007E000FFF0000000FFF;
defparam sdpb_inst_7.INIT_RAM_35 = 256'hF000FFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001F8003FF80;
defparam sdpb_inst_7.INIT_RAM_36 = 256'hFFFFF800FC001FF80000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE003;
defparam sdpb_inst_7.INIT_RAM_37 = 256'hDFEFEFF7FFFFFE003F0007FC00000003FF6FC7EEFFBC1E0F8FE1E0F77C3FBE1F;
defparam sdpb_inst_7.INIT_RAM_38 = 256'hF7BDDFBFD7FBFFFDFFFFFF8007E001FE00000000F7DBEEFB3FEFF7EFDDF77EFE;
defparam sdpb_inst_7.INIT_RAM_39 = 256'hB3EEFF7EFDEFF7FFFDFEFFFFFFFFFFF001F8003F000000003DFBFBBECFBBFDFB;
defparam sdpb_inst_7.INIT_RAM_3A = 256'h03DFCFFDEFF83E1FBF7BEDFFFE7C3FFE1FFFFFFC003F000F800000000F7F7FF7;
defparam sdpb_inst_7.INIT_RAM_3B = 256'h00000000007FF9FF7FFEEFF7FFDEF87F7F5FFFF7FFFFFFFF000FC00000000000;
defparam sdpb_inst_7.INIT_RAM_3C = 256'hF800FE001FFE0000003FFB7FDFBFFFFDFFF7BEFFDFDFFFFDFEFFFFFFE003F000;
defparam sdpb_inst_7.INIT_RAM_3D = 256'hDFEFFFFFFF001F8003FFE000000FFEDFF7DFFFFFFF7EEFBFF7F6FFFF7FBFFFFF;
defparam sdpb_inst_7.INIT_RAM_3E = 256'hBF7EEF0787C3FFFFFFC007E000FFFC000003EF77D9F77FFEDFDFDBEEFDFBBDDF;
defparam sdpb_inst_7.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF000FC003FFF8000007BDFF8FDDFF783F7F1FB;

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[29:0],sdpb_inst_8_dout[1:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_8.READ_MODE = 1'b0;
defparam sdpb_inst_8.BIT_WIDTH_0 = 2;
defparam sdpb_inst_8.BIT_WIDTH_1 = 2;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_8.RESET_MODE = "SYNC";
defparam sdpb_inst_8.INIT_RAM_00 = 256'hFFFFFFE7FFFFE3FE7FFFFFFBFFFFF79FFFFFFFFFE7FFFEFAFFECBFFFF7FEBEFF;
defparam sdpb_inst_8.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF3FFFFF7FD3FFFFF5BFFFFFEAFFFFFFFFFF7FFFFF;
defparam sdpb_inst_8.INIT_RAM_03 = 256'hBFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_04 = 256'hFFAAAEFFB7F7EAEBEBEAFBFBFFFBFFFFFFFFFFFFE1FFFFFDBD7FFFFFCBFFFFFF;
defparam sdpb_inst_8.INIT_RAM_05 = 256'hAFF6BFFFFFBFFFFFF2FFFFFFFFFFFFFFAEFBBFBFBEFFFFFFFFFBDBF5FFFFEFBB;
defparam sdpb_inst_8.INIT_RAM_06 = 256'hFFFFBDEFFFFFFEEBEFFFFFBFFBFFBEFFDBEFEBBE9FFFEFFFFFFFFFFFFF0FFFFD;
defparam sdpb_inst_8.INIT_RAM_07 = 256'hFFFFFFFFFFFE7FFFE4FEFFFFFFCFFFFFFF6FFFFFFFFFF3FFB6EBF6B6F7FBFFBE;
defparam sdpb_inst_8.INIT_RAM_08 = 256'hF2B9A68E34BE7FFA6EA6A7E2FAEBFFEAD6FF3FD8FFCFA7E2EF53AE3FFFFDF9FF;
defparam sdpb_inst_8.INIT_RAM_09 = 256'hAF1EB4F8FE1F800FFFFFFFFFFFFFC2FFFFB3EEFFFFFCBFFFFFD4FFFFFFFFFF7F;
defparam sdpb_inst_8.INIT_RAM_0A = 256'hFFFF2FFFFFFFFFF3FFCF3EEC7FF1DBBF5EFE68774FAC2AFD5DAFF46B245ABC7F;
defparam sdpb_inst_8.INIT_RAM_0B = 256'h98BFFF7EBC677EE3E4C440F383FB39D0FFFFFFFFFFFFFF1FFFFE3FC7FFFFCFFF;
defparam sdpb_inst_8.INIT_RAM_0C = 256'hFFFFD5FDBFFFFD7FFFFFECFFFFFFFFFFFFFB6BE2F7CB7FFFFDAF839B16F116FF;
defparam sdpb_inst_8.INIT_RAM_0D = 256'hFFD8FF7DFCDB274FFF1C7BFB1B7F5EF6FF818F4B771E3BFFFFFFFFFFFFFFFFEE;
defparam sdpb_inst_8.INIT_RAM_0E = 256'h8BDFFFFFFFFFFFFF7FFFFF8BFAFFFFDFFFFFFF8FFFFFFFFFDFFF173F5F3FF2C3;
defparam sdpb_inst_8.INIT_RAM_0F = 256'hEBBFF3A867B3B88FBFF70BF74FC3F7D1FFF4D6FFE3F9FBBFEEEFB0F9F55BCEBD;
defparam sdpb_inst_8.INIT_RAM_10 = 256'hF6BEAB6F0FC57D8ACFBEFFFFFFFFFFFFFEFFFFFDFF93FFFCBFFFFFE0FFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_11 = 256'h9BFFFFFFEFFFFFFFFEFBFEE2AA4BBE1BE5BFEEAB71F4EFF6DFFFAFAFFD27F193;
defparam sdpb_inst_8.INIT_RAM_12 = 256'h1D7FFFFBFFFCFE633F9FFF25F770B7FB0CACBFFFFFFFFFFFFFEFFFFFE3F83FFF;
defparam sdpb_inst_8.INIT_RAM_13 = 256'hFAA9FFFFFE7DFFFFFEFFFFFEBAFFFFFFFF8FFFFCE4F84FE97BA7FEFFB2EF44A8;
defparam sdpb_inst_8.INIT_RAM_14 = 256'hF2B3FF473ABD3957A9DAFFDF9FFFC7FFEFFC66EF96C6613EBCBF0FFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_15 = 256'hCAD2F4BFFFFFFFFBBE5051FFFFF3FBFFFABFFFFFFB9FFFFFFFFCFFFFE317F23B;
defparam sdpb_inst_8.INIT_RAM_16 = 256'hFFFF1BFFFDD6FAB3BFB37D72F0E3FF573E7E3FF5F47FFCBFFCAFDFFEFDF56FF6;
defparam sdpb_inst_8.INIT_RAM_17 = 256'hFECCF33293CC3FDF8F3CBFE6FFFFFFFE80000C2FFFFFC000007FFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_18 = 256'hFFFBFFFFFFFFFFFFFFFFA7FFFFCCCBE1FB24B0BBC34F7DF6BEB1F3FFEADBFFDF;
defparam sdpb_inst_8.INIT_RAM_19 = 256'h17E168FFFDC2FFFDFECA0FDEDA2EEDCCFDEBDCF8FFFFFFFFFFFFFFFDFFFFFCBF;
defparam sdpb_inst_8.INIT_RAM_1A = 256'hFFFFFFFFCFFFFFDFFFFFFFFFFFC5EFFFFFFFF9FFFFFF7F7F75C03F0574FBF2F1;
defparam sdpb_inst_8.INIT_RAM_1B = 256'hFA69A9FFFFBFA0AFF27B6F4EFFBA7FFFCCFBFCE327FE73FCFA483F2FBAFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1C = 256'hFFFEAFFAEFBFFFFFFFFFFFFFFEBFFFFD400002FFFFFA7DFFFFFFE6BBFFFFEC2F;
defparam sdpb_inst_8.INIT_RAM_1D = 256'hFFEA81BFFFFFFFFFBF6FEFFFFEBBF66FEFFF6BBFBFFEFFFFFEAFFFEFAEFFEEFE;
defparam sdpb_inst_8.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAABFFF;
defparam sdpb_inst_8.INIT_RAM_1F = 256'hFFC7FE541D4FF5FDFC55417DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE5FFF;
defparam sdpb_inst_8.INIT_RAM_21 = 256'hFFFFFFFFFFFFF0FFFFFCAA9FFFFF2AAAAAABAAFEAFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFDBFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_26 = 256'hF3FFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFEFFFFEABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFCEFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4FFFFEAFFFFF;
defparam sdpb_inst_8.INIT_RAM_2D = 256'hFFFFFCFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFEBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFFFC7FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7;
defparam sdpb_inst_8.INIT_RAM_34 = 256'hFFFFFFFFFE4FFFFF8BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD8FFFFFDFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_39 = 256'hFFFC2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8BF;
defparam sdpb_inst_8.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFC3FFFFE6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE6FFFFF4FFFFFFFF;

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[29:0],sdpb_inst_9_dout[3:2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_9.READ_MODE = 1'b0;
defparam sdpb_inst_9.BIT_WIDTH_0 = 2;
defparam sdpb_inst_9.BIT_WIDTH_1 = 2;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_9.RESET_MODE = "SYNC";
defparam sdpb_inst_9.INIT_RAM_00 = 256'hFFFFFFF3FFFFFFFEFFFFFFBFFFFFFFCFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF7FFFFF7FEFFFFFFCFFFFFFDFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_03 = 256'h3FFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFF8FF7FFFFFDFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_05 = 256'hFFFFFFFFFDFFFFFFF7FFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFC;
defparam sdpb_inst_9.INIT_RAM_07 = 256'hFFFFFFFFFFFCFFFFF2FFDFFFFFCBFFFFFF3FFFFFFFFFFBFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_08 = 256'hFBFBEFFBEFBEFFFEFFFEBFFFFFABFFEFC7FF802C00E0F7F1EADF2FAFE6F2ABFF;
defparam sdpb_inst_9.INIT_RAM_09 = 256'hAEED3F7A7E9F2AEFFFFFFFFFFFFFF3FFFFFBFCFFFFFF7FFFFFF3FFFFFFFFFFBF;
defparam sdpb_inst_9.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFBDDBEB2ADD7FF6FF9AAFFFFEA3FFE8F3FF2A6CABCAAFF;
defparam sdpb_inst_9.INIT_RAM_0B = 256'hE1F7FF4D7FACD2CBFBE4EDDAFFCFBB31FFFFFFFFFFFFFF0FFFFF7FF3FFFFF7FF;
defparam sdpb_inst_9.INIT_RAM_0C = 256'hFFFFFEFEFFFFFFBFFFFFFEFFFFFFFFFCBFFA73FDD7B1EDFFF3FF494FCEFAB0FF;
defparam sdpb_inst_9.INIT_RAM_0D = 256'hFF8EFEF1FB0FAF2FFC4FFFFF77FF0BEFFFBB9FBF73FEABFF4FFFFFFFFFFFFFF7;
defparam sdpb_inst_9.INIT_RAM_0E = 256'h7DFFFFFFFFFFFFFF2FFFFF1FFBFFFFCBFFFFFFCFFFFFFFFFFFFF1F3F4DFFFFEF;
defparam sdpb_inst_9.INIT_RAM_0F = 256'hFCFFF37BB3D7D9BFFFF1BFFF9F3C7FDBFFEBFEFFF8FFA7BF5FFAF1F0FC8BCFFF;
defparam sdpb_inst_9.INIT_RAM_10 = 256'hFCFFAFBFBFFCBE0FEACFFFFFFFFFFFFFFCFFFFFCFF33FFFEFFFFFFF3FFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_11 = 256'hDFFFFFFF7FFFFFFFFFFFFFF75725FEAEFFFFA2FAECFFD3F2AFFF2F6FFFBBF6B7;
defparam sdpb_inst_9.INIT_RAM_12 = 256'hFEFFF2FEFFFCFF96BFDFF63DF6FE33F3FD01FFFFFFFFFFFFFFDFFFFFFFF33FFF;
defparam sdpb_inst_9.INIT_RAM_13 = 256'hFFFE3FFFFFFFBFFFFEFFFFFFF7FFFFFFFFF7FFFDB8BEDFCA5F0FFFEFEEBFB5EF;
defparam sdpb_inst_9.INIT_RAM_14 = 256'hF5F5DB99FC7E739EE9FBFF8FFFFFDFFFFBFDFFFBF3A78A3E42BFB7FFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_15 = 256'hDFC3F4BFFFFFFFFD4557F7FFFFF90FFFFFBFFFFFFCCFFFFFFFFCFFFFDFF3D4BF;
defparam sdpb_inst_9.INIT_RAM_16 = 256'hFFFF7FFFFEEFFE13FF7F3FF7ADD7EBBAFD7D7FFF76FFFCFFFCAFF7FE7EBD3A37;
defparam sdpb_inst_9.INIT_RAM_17 = 256'hF56BF93173F3D3BFCE7C3FC7FFFFFFFFC7FFF7FFFFFFFFFFFFF7FFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_18 = 256'hFFFFFFFFFFFBFFFFFFFFF7FFFFDBA3FF7E03BABF4E3C3C33FBFBEBFFE82FFFEE;
defparam sdpb_inst_9.INIT_RAM_19 = 256'hA7FBABBFFCEEFFFDEF7FFFF77F3DE9F8F0D7EFFAFFFFFFFFFFFFFFFDFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_1A = 256'hFFFFFFFFEFFFFFFFFFFFFFFFFFE63FFFFFFFFDFFFFFF6ABF53DAAB8BF6F6EFCF;
defparam sdpb_inst_9.INIT_RAM_1B = 256'hFEFFFE7DAFDFFEFDFBFC3E1FFFF43FFFF3F803FCFC03FCBF2F7EBF7FDBFFFFFF;
defparam sdpb_inst_9.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC6AAAAA55555FFCFFFFFFFE3FFFFFFD4F;
defparam sdpb_inst_9.INIT_RAM_1D = 256'hFFFFFDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_1F = 256'hFFE3FF000C0FF0FCFC0019BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFF;
defparam sdpb_inst_9.INIT_RAM_21 = 256'hFFFFFFFFFFFFFCFFFFFCA5500000555556A9AAFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCCFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDCFFFFCFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_26 = 256'hFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFBFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFCEFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFCFFFFF;
defparam sdpb_inst_9.INIT_RAM_2D = 256'hFFFFFDFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFF3FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFF;
defparam sdpb_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFF7FFFFF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFCFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_39 = 256'hFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3F;
defparam sdpb_inst_9.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFF7FFFFFFFF;

SDPB sdpb_inst_10 (
    .DO({sdpb_inst_10_dout_w[29:0],sdpb_inst_10_dout[5:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_10.READ_MODE = 1'b0;
defparam sdpb_inst_10.BIT_WIDTH_0 = 2;
defparam sdpb_inst_10.BIT_WIDTH_1 = 2;
defparam sdpb_inst_10.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_10.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_10.RESET_MODE = "SYNC";
defparam sdpb_inst_10.INIT_RAM_00 = 256'hFFFFFFF2AAAAA7FDAAAAAAFFFFFFFABAAAAAAAAAA3FFFFFFFFFFBFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF2AAAAA7FFEAAAAAAFFFFFFCAAAAAAAAAAA7FFFFF;
defparam sdpb_inst_10.INIT_RAM_03 = 256'h2AAAAAAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBAAAAABFF6AAAAABFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_05 = 256'hBFF2AAAAA8FFFFFFFAAAAAAAAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCAAAAB;
defparam sdpb_inst_10.INIT_RAM_07 = 256'hFFFFFFFFFFFCAAAAADFFFAAAAABFFFFFFF6AAAAAAAAAA3FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF5FFFFBFFFFFFFFFFFFAFFFFBFBEFEFFBFEABFF;
defparam sdpb_inst_10.INIT_RAM_09 = 256'h6E9DFAF2FDBF2AFFFFFFFFFFFFFFFEAAAAAFFFAAAAAAFFFFFFFEAAAAAAAAAA7F;
defparam sdpb_inst_10.INIT_RAM_0A = 256'hFFFFEAAAAAAAAAABFFBFFC7D3AABFFFF6FFBA8FEBFEA2FFDBD7FF2AACA8CAA7F;
defparam sdpb_inst_10.INIT_RAM_0B = 256'hEEC3FFA3BFA4E9ABFFFCFBD96BDAFAEFFFFFFFFFFFFFFFBAAAAAFFDEAAAAAFFF;
defparam sdpb_inst_10.INIT_RAM_0C = 256'hAAAAAFFFAAAAAAFFFFFFFFAAAAAAAAABFFF3FDEBD719AE7FF6FF36FFF8FF52FF;
defparam sdpb_inst_10.INIT_RAM_0D = 256'hFF3DF2F6FE5FC34FFFDEBFFF7FFFFFFBFF2FFFDFEA7CF3FFEFFFFFFFFFFFFFF2;
defparam sdpb_inst_10.INIT_RAM_0E = 256'hF0FFFFFFFFFFFFFFEAAAAAEFFAAAAABFFFFFFFFAAAAAAAAAAFFFBB7F0DBFE9C3;
defparam sdpb_inst_10.INIT_RAM_0F = 256'hABFFFEBAF8DFFF8EBFF35F6BDFE3FFF7FFFFFAFFFBBFAABFEFF6BAF4FD33CE7F;
defparam sdpb_inst_10.INIT_RAM_10 = 256'hF0FFA70F8FEBFF3BCAAFFFFFFFFFFFFFFEAAAAABFFAEAAA8FFFFFFFEAAAAAAAA;
defparam sdpb_inst_10.INIT_RAM_11 = 256'h8FFFFFFF2AAAAAAAAA3FFFE7FBBDFFABFAFFFBFF24FA53FE8FFF6F0FFFEBF2A7;
defparam sdpb_inst_10.INIT_RAM_12 = 256'hA6FFFDF6FFFC3F3CBF6FFE7BFFFC2BE37EA4FFFFFFFFFFFFFFEAAAAAAFFAEAAA;
defparam sdpb_inst_10.INIT_RAM_13 = 256'hFFFF2AAAAA3F6AAAABFFFFFFF6AAAAAAAAA3FFFDFC3C53CA2F1FF8C7DAAFA9BC;
defparam sdpb_inst_10.INIT_RAM_14 = 256'hF4F7EBB8FE2BBA59FEFFFF4FBFFFEBFFFFF8FFEFEF3FF37ED3FF6FFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_15 = 256'hEABBFBBFFFFFFFFF5003FEAAAAAC5AAAAA7FFFFFFEBAAAAAAAA9FFFFF7CFC57F;
defparam sdpb_inst_10.INIT_RAM_16 = 256'hAAAAEFFFFDBC7EFBFFEF8C3AAAF7C36AAD3FFFFEBFFFFC3FFDBFFFFEBCF3F2EF;
defparam sdpb_inst_10.INIT_RAM_17 = 256'hFC0AF7F037EF3FCFBDBDFFB7FFFFFFFFEFFFFFEAAAAABFFFFFDFFFFFFFAAAAAA;
defparam sdpb_inst_10.INIT_RAM_18 = 256'hFFFFFFFFFFE2AAAAAAAAA7FFFFFD3BFEBCAABF7F7FFD3EB6B6FE3FFFDC3FFFDB;
defparam sdpb_inst_10.INIT_RAM_19 = 256'h2FF32A7FFEA8FFFEAFEA9FAB6AFF2AE8F1DFDBFFFFFFFFFFFFFFFFFCAAAAAAFF;
defparam sdpb_inst_10.INIT_RAM_1A = 256'hFFFFFFFFFAAAAA8FFFFFFFFFFFF3EAAAAAAAA9FFFFFF2A7F6FDAA3CA73F3DBFF;
defparam sdpb_inst_10.INIT_RAM_1B = 256'hFEFFAAFF1FBFEFBFBEFFFE6FFFFDBFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFDAAAAABAAAAA800000EABAAAAAAA8FFFFFFFE2F;
defparam sdpb_inst_10.INIT_RAM_1D = 256'hAAAAA97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_10.INIT_RAM_1F = 256'hAABEAAFFFBFAAFABABFFF4BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2AAA;
defparam sdpb_inst_10.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDBAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBAAAA9FFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_26 = 256'hEAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFF6AAAAA3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7AAAABBFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBAAAAAAFFFFF;
defparam sdpb_inst_10.INIT_RAM_2D = 256'hFFFFFCAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFDAAAAA8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2AAAAABFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAA7;
defparam sdpb_inst_10.INIT_RAM_34 = 256'hFFFFFFFFFF6AAAAA3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_39 = 256'hAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEA;
defparam sdpb_inst_10.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFEAAAAA3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAABFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAFFFFFFFFF;

SDPB sdpb_inst_11 (
    .DO({sdpb_inst_11_dout_w[29:0],sdpb_inst_11_dout[7:6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_11.READ_MODE = 1'b0;
defparam sdpb_inst_11.BIT_WIDTH_0 = 2;
defparam sdpb_inst_11.BIT_WIDTH_1 = 2;
defparam sdpb_inst_11.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_11.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_11.RESET_MODE = "SYNC";
defparam sdpb_inst_11.INIT_RAM_00 = 256'hFFFFFFF955555FFF5555557FFFFFFD55555555555BFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFD55555BFF5555557FFFFFFF55555555555BFFFFF;
defparam sdpb_inst_11.INIT_RAM_03 = 256'h95555555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555557FF9555556FFFFFFF;
defparam sdpb_inst_11.INIT_RAM_05 = 256'h6FFD555556FFFFFFF95555555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE55555;
defparam sdpb_inst_11.INIT_RAM_07 = 256'hFFFFFFFFFFFF555556FFD555555FFFFFFFD5555555555FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_09 = 256'hAF7F7DBDFF6FD57FFFFFFFFFFFFFF555555FFE555555FFFFFFFD5555555555FF;
defparam sdpb_inst_11.INIT_RAM_0A = 256'hFFFFD5555555555FFF9F6EBEB957DBFFDBFD57FD7FE5BFFF7EBFFD56E56F55BF;
defparam sdpb_inst_11.INIT_RAM_0B = 256'hF7FBFFE9AEAAFA6BF9F7F7F7DFF5FEA7FFFFFFFFFFFFFF955555BFF555555FFF;
defparam sdpb_inst_11.INIT_RAM_0C = 256'h555557FF555555FFFFFFFD5555555555FFFDFAF7EBEA7EBFFD7FDA6FD7FDBAFF;
defparam sdpb_inst_11.INIT_RAM_0D = 256'hFFD7FDFAFDAFEFEFFF7F7FFFDFFFDFF7FFDF6F7F9DFF5FFF7FFFFFFFFFFFFFFD;
defparam sdpb_inst_11.INIT_RAM_0E = 256'hFBFFFFFFFFFFFFFFD555557FF955555FFFFFFFD5555555556FFFDFDFBEBFF7FB;
defparam sdpb_inst_11.INIT_RAM_0F = 256'h57FFFDFDFAEBFF7F7FFDAFDFAFDDFFF9FFF6F7FFFDFFFDFF7FFDFAFBFE9FF6BF;
defparam sdpb_inst_11.INIT_RAM_10 = 256'hFBFFDFEFAFE5BEB7F56FFFFFFFFFFFFFFE555556FFD55556FFFFFFFD55555555;
defparam sdpb_inst_11.INIT_RAM_11 = 256'h7FFFFFFFD555555555BFFFDFDFDEBD56F7FF9DFDAAFDEFF96FFFAFBFFFDFF95F;
defparam sdpb_inst_11.INIT_RAM_12 = 256'h5BFFFAFAFFFEFFEABFAFFDFDF9FE9BEBAFAAFFFFFFFFFFFFFFF555555FFD5555;
defparam sdpb_inst_11.INIT_RAM_13 = 256'hFFFF955555FF955557FFFFFFF9555555555FFFFEBEFEEFFAAFBFFAEFF55FDF7F;
defparam sdpb_inst_11.INIT_RAM_14 = 256'hFEFAEF9A7EBDFDA7E7FFFFEF9FFFEBFFE7FAFFDBDFDFDEBE69FFDFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_15 = 256'hE55FFDFFFFFFFFFEAAA955555556A55555BFFFFFFF5555555556FFFFEBEBFAFF;
defparam sdpb_inst_11.INIT_RAM_16 = 256'h55557FFFFF7EBF5FFFDFAEF957EBEFD56FBE7FFDF9FFFFBFFF7F9FFEBEBDFDF7;
defparam sdpb_inst_11.INIT_RAM_17 = 256'hFAA7FDFE9BE69F6F7EBEBFDFFFFFFFFFE555555555555555556FFFFFFFD55555;
defparam sdpb_inst_11.INIT_RAM_18 = 256'hFFFFFFFFFFF9555555555FFFFFF6DBF5FFA9F9DBAF6FBEBDFDF6D7FFE79FFFF7;
defparam sdpb_inst_11.INIT_RAM_19 = 256'hDFDFD5FFFF57FFFF7F957FDFD57F96F7FBEBF7FDBFFFFFFFFFFFFFFE555557FF;
defparam sdpb_inst_11.INIT_RAM_1A = 256'hFFFFFFFFE555556FFFFFFFFFFFFD5555555557FFFFFFD5FFDFF55FE5FAFDF7E7;
defparam sdpb_inst_11.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF555555AAAAAAAAAAA55555555556FFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1D = 256'h555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF555555555555555555555;
defparam sdpb_inst_11.INIT_RAM_1F = 256'h555555555555555555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555;
defparam sdpb_inst_11.INIT_RAM_21 = 256'hFFFFFFFFFFFFFD555557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE555556FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE555556FFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_26 = 256'hF555555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFF955555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555557FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555557FFFFF;
defparam sdpb_inst_11.INIT_RAM_2D = 256'hFFFFFE555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFF555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF955555FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF955555B;
defparam sdpb_inst_11.INIT_RAM_34 = 256'hFFFFFFFFFFD55555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFD555557FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE555556FFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_39 = 256'h5555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF55;
defparam sdpb_inst_11.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFF555555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF955555BFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD555557FFFFFFFF;

SDPB sdpb_inst_12 (
    .DO({sdpb_inst_12_dout_w[27:0],sdpb_inst_12_dout[3:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_12.READ_MODE = 1'b0;
defparam sdpb_inst_12.BIT_WIDTH_0 = 4;
defparam sdpb_inst_12.BIT_WIDTH_1 = 4;
defparam sdpb_inst_12.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_12.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_12.RESET_MODE = "SYNC";
defparam sdpb_inst_12.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_01 = 256'hFFFFF1FFFFFFFFFFE2FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7EFFFFFFFFFF4CEFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_08 = 256'hFFFFFFFFF7CFFFFFFFFFF6DEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFEBFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_0F = 256'hFFFFFFFFFFFFFF6DFFFFFFFFFF2EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2A0FFFFFFFFFC1FF;
defparam sdpb_inst_12.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFECEFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_19 = 256'hEDFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1DFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_20 = 256'hFFFF0F5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFF;
defparam sdpb_inst_12.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDFCFFFFFFFFFF67FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_27 = 256'hFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE4;
defparam sdpb_inst_12.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE3D0EFFFFFFFFDFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2E = 256'hFFFCAF1FFFFFFFFECFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE4DEFFFFFFFFF9FFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_35 = 256'hFFFFFFFFF7FFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0EFFFFFFFFFEFEFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3C = 256'hFFFFFFFFFFFFFBFFFFFFFFFFE2EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_13 (
    .DO({sdpb_inst_13_dout_w[27:0],sdpb_inst_13_dout[7:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_13.READ_MODE = 1'b0;
defparam sdpb_inst_13.BIT_WIDTH_0 = 4;
defparam sdpb_inst_13.BIT_WIDTH_1 = 4;
defparam sdpb_inst_13.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_13.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_13.RESET_MODE = "SYNC";
defparam sdpb_inst_13.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_01 = 256'hFFFFF966666666666CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB666666666668FFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_08 = 256'hFFFFFFFFFE666666666667EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF866666666666CFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFD666666666668FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF776666666666EFF;
defparam sdpb_inst_13.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFF866666666666AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_19 = 256'h68FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD6666666666;
defparam sdpb_inst_13.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFF766666666666EFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_20 = 256'h666676AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB66666;
defparam sdpb_inst_13.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFD666666666667FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_27 = 256'h66666666667DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam sdpb_inst_13.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE67666666666AFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2E = 256'hFFFF867666666666FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC66666666666CFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_35 = 256'hFFFFFFFFF866666666669FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD66666666667FFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3C = 256'hFFFFFFFFFFFFFF76666666666DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_14 (
    .DO({sdpb_inst_14_dout_w[23:0],sdpb_inst_14_dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_1}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_14.READ_MODE = 1'b0;
defparam sdpb_inst_14.BIT_WIDTH_0 = 8;
defparam sdpb_inst_14.BIT_WIDTH_1 = 8;
defparam sdpb_inst_14.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_14.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_14.RESET_MODE = "SYNC";
defparam sdpb_inst_14.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE736F6E6F6F6F6F6F6F6F87FFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAB6C716F6F6F6F6F6F6F6CEAFF;
defparam sdpb_inst_14.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0D = 256'hC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFE896E6F6F6F6F6F6F6F6F;
defparam sdpb_inst_14.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_14 = 256'h6F6F93FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC746E6E6F6F6F6F;
defparam sdpb_inst_14.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1B = 256'h6F6F6F6E6CEEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE4736E6F6F;
defparam sdpb_inst_14.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_22 = 256'h6E6F6F6F6F6F6EB2FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFD76D;
defparam sdpb_inst_14.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_29 = 256'hFEEB7C6C6F6E6F6F6F88FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_30 = 256'hFFFFFEFEFCB96F6B6D6E6E6EF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_37 = 256'hFFFFFFFFFEFFFEFFF8D5BE9CA2BBEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_14.INIT_RAM_3D = 256'h00000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sdpb_inst_12_dout[0]),
  .I1(sdpb_inst_14_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(sdpb_inst_8_dout[0]),
  .I1(mux_o_6),
  .S0(dff_q_1)
);
MUX2 mux_inst_9 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(mux_o_8),
  .S0(dff_q_0)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(sdpb_inst_12_dout[1]),
  .I1(sdpb_inst_14_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(sdpb_inst_8_dout[1]),
  .I1(mux_o_16),
  .S0(dff_q_1)
);
MUX2 mux_inst_19 (
  .O(dout[1]),
  .I0(sdpb_inst_1_dout[1]),
  .I1(mux_o_18),
  .S0(dff_q_0)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(sdpb_inst_12_dout[2]),
  .I1(sdpb_inst_14_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(sdpb_inst_9_dout[2]),
  .I1(mux_o_26),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(dout[2]),
  .I0(sdpb_inst_2_dout[2]),
  .I1(mux_o_28),
  .S0(dff_q_0)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(sdpb_inst_12_dout[3]),
  .I1(sdpb_inst_14_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(sdpb_inst_9_dout[3]),
  .I1(mux_o_36),
  .S0(dff_q_1)
);
MUX2 mux_inst_39 (
  .O(dout[3]),
  .I0(sdpb_inst_3_dout[3]),
  .I1(mux_o_38),
  .S0(dff_q_0)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sdpb_inst_13_dout[4]),
  .I1(sdpb_inst_14_dout[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(sdpb_inst_10_dout[4]),
  .I1(mux_o_46),
  .S0(dff_q_1)
);
MUX2 mux_inst_49 (
  .O(dout[4]),
  .I0(sdpb_inst_4_dout[4]),
  .I1(mux_o_48),
  .S0(dff_q_0)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(sdpb_inst_13_dout[5]),
  .I1(sdpb_inst_14_dout[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(sdpb_inst_10_dout[5]),
  .I1(mux_o_56),
  .S0(dff_q_1)
);
MUX2 mux_inst_59 (
  .O(dout[5]),
  .I0(sdpb_inst_5_dout[5]),
  .I1(mux_o_58),
  .S0(dff_q_0)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(sdpb_inst_13_dout[6]),
  .I1(sdpb_inst_14_dout[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(sdpb_inst_11_dout[6]),
  .I1(mux_o_66),
  .S0(dff_q_1)
);
MUX2 mux_inst_69 (
  .O(dout[6]),
  .I0(sdpb_inst_6_dout[6]),
  .I1(mux_o_68),
  .S0(dff_q_0)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(sdpb_inst_13_dout[7]),
  .I1(sdpb_inst_14_dout[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(sdpb_inst_11_dout[7]),
  .I1(mux_o_76),
  .S0(dff_q_1)
);
MUX2 mux_inst_79 (
  .O(dout[7]),
  .I0(sdpb_inst_7_dout[7]),
  .I1(mux_o_78),
  .S0(dff_q_0)
);
endmodule //Gowin_SDPB1
