//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Sun Aug 06 14:52:33 2023

module Gowin_pROM1 (dout, clk, oce, ce, reset, ad);//grayscale etf

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [16:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [1:1] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [1:1] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [1:1] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [1:1] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [2:2] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [2:2] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [2:2] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [2:2] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [3:3] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [3:3] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [3:3] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [3:3] prom_inst_15_dout;
wire [30:0] prom_inst_16_dout_w;
wire [0:0] prom_inst_16_dout;
wire [30:0] prom_inst_17_dout_w;
wire [1:1] prom_inst_17_dout;
wire [30:0] prom_inst_18_dout_w;
wire [2:2] prom_inst_18_dout;
wire [30:0] prom_inst_19_dout_w;
wire [3:3] prom_inst_19_dout;
wire [29:0] prom_inst_20_dout_w;
wire [1:0] prom_inst_20_dout;
wire [29:0] prom_inst_21_dout_w;
wire [3:2] prom_inst_21_dout;
wire [27:0] prom_inst_22_dout_w;
wire [3:0] prom_inst_22_dout;
wire [30:0] prom_inst_23_dout_w;
wire [4:4] prom_inst_23_dout;
wire [30:0] prom_inst_24_dout_w;
wire [4:4] prom_inst_24_dout;
wire [30:0] prom_inst_25_dout_w;
wire [4:4] prom_inst_25_dout;
wire [30:0] prom_inst_26_dout_w;
wire [4:4] prom_inst_26_dout;
wire [30:0] prom_inst_27_dout_w;
wire [5:5] prom_inst_27_dout;
wire [30:0] prom_inst_28_dout_w;
wire [5:5] prom_inst_28_dout;
wire [30:0] prom_inst_29_dout_w;
wire [5:5] prom_inst_29_dout;
wire [30:0] prom_inst_30_dout_w;
wire [5:5] prom_inst_30_dout;
wire [30:0] prom_inst_31_dout_w;
wire [6:6] prom_inst_31_dout;
wire [30:0] prom_inst_32_dout_w;
wire [6:6] prom_inst_32_dout;
wire [30:0] prom_inst_33_dout_w;
wire [6:6] prom_inst_33_dout;
wire [30:0] prom_inst_34_dout_w;
wire [6:6] prom_inst_34_dout;
wire [30:0] prom_inst_35_dout_w;
wire [7:7] prom_inst_35_dout;
wire [30:0] prom_inst_36_dout_w;
wire [7:7] prom_inst_36_dout;
wire [30:0] prom_inst_37_dout_w;
wire [7:7] prom_inst_37_dout;
wire [30:0] prom_inst_38_dout_w;
wire [7:7] prom_inst_38_dout;
wire [30:0] prom_inst_39_dout_w;
wire [4:4] prom_inst_39_dout;
wire [30:0] prom_inst_40_dout_w;
wire [5:5] prom_inst_40_dout;
wire [30:0] prom_inst_41_dout_w;
wire [6:6] prom_inst_41_dout;
wire [30:0] prom_inst_42_dout_w;
wire [7:7] prom_inst_42_dout;
wire [29:0] prom_inst_43_dout_w;
wire [5:4] prom_inst_43_dout;
wire [29:0] prom_inst_44_dout_w;
wire [7:6] prom_inst_44_dout;
wire [27:0] prom_inst_45_dout_w;
wire [7:4] prom_inst_45_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire dff_q_6;
wire dff_q_7;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_88;
wire mux_o_89;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_0.INIT = 16'h0002;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_1.INIT = 16'h0008;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_2.INIT = 16'h0020;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_3.INIT = 16'h0080;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_4.INIT = 16'h0200;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad[13]),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16])
);
defparam lut_inst_5.INIT = 16'h0400;
LUT2 lut_inst_6 (
  .F(lut_f_6),
  .I0(ce),
  .I1(lut_f_5)
);
defparam lut_inst_6.INIT = 4'h8;
LUT5 lut_inst_7 (
  .F(lut_f_7),
  .I0(ad[12]),
  .I1(ad[13]),
  .I2(ad[14]),
  .I3(ad[15]),
  .I4(ad[16])
);
defparam lut_inst_7.INIT = 32'h00400000;
LUT2 lut_inst_8 (
  .F(lut_f_8),
  .I0(ce),
  .I1(lut_f_7)
);
defparam lut_inst_8.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b1;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE5F93BFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFE;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDDB2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7F3FBF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF3FF4C7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FF8FFFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFBFFF8B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3FFFE7FFFFFF;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFF6FFFEB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDBFFF91FFFFFFFFF;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFF3FFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFF1FFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFEFFFFDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFA77FFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFF9FFFD0BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFF473FFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFFFFFEFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE6FFFF0BFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFEBFFFF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE5FFFF8F3FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1E = 256'hFC7FFFF48FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE17FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFFABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFB3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFEDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE3FFFFA7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE6FFFFE9FFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFF97FFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFEFFFFFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFF9FFFFFFFFF;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFF9FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFF9FFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFF27FFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCDFFFFC7FFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFFFFFF27FFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC9FFFFEBFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFF07FFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC2FFFFC33FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFF2FFFFFF4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b1;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFE4FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hEBFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFFF33FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDF;
defparam prom_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFDDFFFFB7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_07 = 256'hFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFDF;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFF7FFF;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFC7FFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFF77FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFEBFFFFBCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFE43FFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFEBFFFFC5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFFEBFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFFFFBFFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFDFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFFEFFFFEAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF86FFFFFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hFFEFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5FFFFDFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_24 = 256'hFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFF0BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCBF;
defparam prom_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFD0FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFF;
defparam prom_inst_1.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFF8FFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFFFFFDC67CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFF6FFFFE3F;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFEFFFFFFFFFFFFCBFFFFFFFFFFFE39E2EFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_30 = 256'h0143F3AE8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF60000000000004FFFFFC0000;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFB7FFFFFFFFFFFE7FFFFC7FFFFF57C1E243FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFD9E67FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hBFFFFFFFFFFFFFFAFFFFFFCEFFFB7B27EFFFEC3FFFFFFFFFFFFFFFFFE7FFFC7B;
defparam prom_inst_1.INIT_RAM_35 = 256'h9FFE2000000000000BFFFFF40000E1FFFF820403FFFFFEE7FFFFFFFFFF9FFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hFF077E3FFFF81B7A8369FFCFEBDF4D96DF9F7F01C84625822F3D0205E5C33D85;
defparam prom_inst_1.INIT_RAM_37 = 256'hF3BFF04A0108C8DB1D52D3E331A60E57FEB80000000000017FFFFE00015FFFFF;
defparam prom_inst_1.INIT_RAM_38 = 256'hEA7FFFFFFFFFFF3FFFFF8FFFF5FFFFFFFF18CFFFFEC25E30033FF3F8D1EBFC37;
defparam prom_inst_1.INIT_RAM_39 = 256'hE73FFFFF03B1D30A87F87EAA70FF99FDFDD6B701C30230C8564ABC29194FAEFF;
defparam prom_inst_1.INIT_RAM_3A = 256'hFC297F71F8E6D56BAB9FA923FCB3FFF180000000000017FFFFCE001EBFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'h000000000007FFFFF0000677FFFFFFFDCFFBFFE87CF6BDB5FDBFFEDD6FD9FEFB;
defparam prom_inst_1.INIT_RAM_3C = 256'h357FFC177901A4FF63C827378EBFCF9B7140DEF413D0771F8FF349F11F2FFFD8;
defparam prom_inst_1.INIT_RAM_3D = 256'hDBE5E94C7AE1AFA6DFCD3C5EDBFFEFFFFFFFFFFFFE5FFFFC0000CC9FFFFFFFF9;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFFFFFC7FFFFFFFFFCFFFFFFFFFE49BFFFDFEAD7D0F7C0138BFDFBC7F7CEFD;
defparam prom_inst_1.INIT_RAM_3F = 256'hFF16BBB7F177FB2678F5FE73FAF5FF3FF3E15FBF9E4BE2B779DF9D9CFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b1;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hF19E46F711FA69FD59679ABFFFFFFFFFFFFFFFFCFFFFE9FFFC87FFFFFFFF967F;
defparam prom_inst_2.INIT_RAM_01 = 256'hFFFFFC7FFFFCFFFFC6FFFFFFFFFE1FFFDFCF3DFFFEFC61EBFFCE7EFF9C5FCBFF;
defparam prom_inst_2.INIT_RAM_02 = 256'hE51F7F577F3FD7B7DFA7FFBE57F0FFDEF515B9403A9A77BB4C88FFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_03 = 256'hD732F64801C8ECF973A97FFE0000001800BFFFFFFE5FFFF59FFFFFFFFF84FFFE;
defparam prom_inst_2.INIT_RAM_04 = 256'hABE3FFFFCFFFFFA6FFFFFFFFF8BFFF7CBBFE977FC23A2FFECB0FFB93FC3F139D;
defparam prom_inst_2.INIT_RAM_05 = 256'h37EDF7F30DEA7C8C13FCEBFF28E0CE7FC7764E04BE34955EEA1FFFCC00080E03;
defparam prom_inst_2.INIT_RAM_06 = 256'h7CD0823BAEF837BF43FFF0FFFBFFFFAA7E3FFFFD7FFFF83FFFFFFFFFE7FFB709;
defparam prom_inst_2.INIT_RAM_07 = 256'h5BFFFE7FFFFF9FFFFFFFFFE3FFFDF169D9F9FDE8113F509BFF13BFEE7030BE7E;
defparam prom_inst_2.INIT_RAM_08 = 256'h3AFF71080DBCA2BFD3CBF8B465B7BE1F71E022BB3FC55FDCFFFF00015F9FF51E;
defparam prom_inst_2.INIT_RAM_09 = 256'h6A375686B2B8F3BFFF7FFFAFFFFEC3ABFFFF87FFFFD7FFFFFFFFF07FFEFDFF70;
defparam prom_inst_2.INIT_RAM_0A = 256'hFFFDFFFFF7FFFFFFFFFE9FFF3DEAB98213D660BDFFCC7FFF7AFFAAA207F39AEF;
defparam prom_inst_2.INIT_RAM_0B = 256'hF01F9FFFCF5C7FC93F07FDF2FFF5FEC579713C695C4EAFFFBFFFFBFF03C4EF7F;
defparam prom_inst_2.INIT_RAM_0C = 256'h91CE4117982FFFFFFFF9FFFFF9FFDFFFFC1FFFFDBFFFFFFFFF6DFFC7BF7E7E03;
defparam prom_inst_2.INIT_RAM_0D = 256'h31FFFFEFFFFFFFFFFFFFFCB2DFFFA27DA22EEB25839E73DFC9BEC2BE9E13B3BC;
defparam prom_inst_2.INIT_RAM_0E = 256'hA4A6E21AEB9CDFF87F85FBDDE38F6F657B222DA537FFFFFFFFCFFFFF5FC7FFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'hDD12D76AFFFFFFFF87FFFFFFF7FFFFCCFFFFEDFFFFFFFFFEA3FD8DBC7FFF387A;
defparam prom_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFA9FF21713FFECA16557858BD74F978FE9FF977E7F83E6EEBE4;
defparam prom_inst_2.INIT_RAM_11 = 256'h71CC5BBF3FBF8FD88F39BF03D030E0A148A7C53FFFFFFFECBFFFF5FEBFFFFA3F;
defparam prom_inst_2.INIT_RAM_12 = 256'h3DFA2FFFFFFFFB47FFFF77CFFFFFAFFFFFFFFFFFFFFFEE7FEEB4B7FECBA07F24;
defparam prom_inst_2.INIT_RAM_13 = 256'hE7FFFFFFFFFF0FFE8EB9FFD0901C4D7573652FDE2FC9F4AF4E73DC45EC33C9EF;
defparam prom_inst_2.INIT_RAM_14 = 256'h03B7FABBF1BC75CFA2091A6C0363EB6FB9E5FFFFFFFFFEFFFFBFE7FFFFCDFFFF;
defparam prom_inst_2.INIT_RAM_15 = 256'hC7FFFFFFFFFE3FFFE0EE3FFFF3FFFFFFFFFFFFFFFFDCFE881BBEFA6C4735D57D;
defparam prom_inst_2.INIT_RAM_16 = 256'hFFFFFFFFFADFD2565F9FF0F3EDEEF7F3F5FFFCFFEF2EF4FDC08C8F5AE3F053AE;
defparam prom_inst_2.INIT_RAM_17 = 256'h3F47FFE7D83E5AC78AADA8381D2B7460DFFFFFFFFFC7FFFDF89FFFFF7FFFFFFF;
defparam prom_inst_2.INIT_RAM_18 = 256'hFFFFFFFFFFFFFE7E17FFFFAFFFFFBFFFFFFFFFFEDFF0499408612A7D13CBF914;
defparam prom_inst_2.INIT_RAM_19 = 256'hFFFFFF5FFDE8600FF0B79F4AF37F056FFB9FFC77FF2AA3E67AC3C647F31F0C87;
defparam prom_inst_2.INIT_RAM_1A = 256'hFFFE3C7FD47C79ACA2EDB9FE9FF50FFFFFFFFFE6FFFF8FF0FFFFFA7FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1B = 256'hFFFFFF6FFFF0FBFFFFFC9FFFF7FFFFFFFFFFF9FF743D03ECC2239EBD9DE013F0;
defparam prom_inst_2.INIT_RAM_1C = 256'hFFFFDFFFBFF2F7037DEFFF77FE17FC79FFD7FFFAFFFEEFFE3CFF7F7FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDFFFEBFCFFFFFA3FFFD7FFFFFFF;
defparam prom_inst_2.INIT_RAM_1E = 256'hFFFBFFFF9FE1FFFFEDFFFEBFFFFFFFFFFFE7FFFFFFFD4BFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1F = 256'hF3FFFFFFFF403FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF85FFFFBFFFFFFF87FFFDFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_21 = 256'hEFFFFC7EBFFFFE1FFFABFFFFFFFFFFFCCFFFFFFFF20FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_22 = 256'hF9EF3E71EFEFA7FEFFFFFFFCFF9FFFCFBFFFFFF1FEFFFFFFF33FFF3FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_23 = 256'h4FDC003FCFE83FFD2F506FFFFFFFFFFCFFFF5FC3FFFFEFFFEAFFFFFFFFFFFF13;
defparam prom_inst_2.INIT_RAM_24 = 256'hFFE3F9FFFFFDFFF55FFFFFFFFFFFF3E6618C9C899B7A3FDFCFF00F01D79DB3E4;
defparam prom_inst_2.INIT_RAM_25 = 256'h3D3F53CEE5C7E72FEC0FE80EE20DFB13FA029281F60BFF87C817FFFFFFFFFC7F;
defparam prom_inst_2.INIT_RAM_26 = 256'h80A4A9FE06EFF6F71BFFFFFFFFFFDFFFF8BC3FFFFE7FFF7FFFFFFFFFFFFAB0F6;
defparam prom_inst_2.INIT_RAM_27 = 256'h9D97FFFFFFFF5BFFFFFFFFFFFEADBEBFDFCED99403FDD0F9037C3F7A8B7F82BF;
defparam prom_inst_2.INIT_RAM_28 = 256'h734475F07E743F7FBF609ED36FF73F70A0873F9E37EFBE7EFFFFFFFFFFEFFFFC;
defparam prom_inst_2.INIT_RAM_29 = 256'hC5BFEF2EF8FFAF2FFFFFFFFFFDFFFF4319FFFFDA67FDFFFFFFFFFFFFA6C39781;
defparam prom_inst_2.INIT_RAM_2A = 256'hFFFFF218477FFFFFFFFFFFFFFAFC435CE03CAB579537CF078FB7DB37D445FB32;
defparam prom_inst_2.INIT_RAM_2B = 256'h0E6B6FED55F58BE171ED74F4767517E69EF629FEAFF723FFFFFFFFFFDFFFFDC5;
defparam prom_inst_2.INIT_RAM_2C = 256'h5C76BFADF9D9FFFFFFFFFF87FFFDEB6FFFFF072BFFFFFFFFFFFFFEFCFEDBFFAE;
defparam prom_inst_2.INIT_RAM_2D = 256'hFFD7F33FFFFFFFFFFFFFEF0FCB65E013FFABFDDFFFE57FB9FFFD3D920DAD3E1F;
defparam prom_inst_2.INIT_RAM_2E = 256'h955E5F7FDC3FF9FF391FFFF3FE7F126F5EFFFF3FFF3FFFFFFFFFF8FFFF3BD7FF;
defparam prom_inst_2.INIT_RAM_2F = 256'hD3FFEFEF8FFFFFFFFFFC7FFFFAF17FFFFEFDEFFFFFFFFFFFFFE7DBFE9D7878FC;
defparam prom_inst_2.INIT_RAM_30 = 256'hF8EBFFFFFFFFFFFFFDF0FE115EDADD7CB7B38FFE6FF83FED4FE8CFFF5FECCFE3;
defparam prom_inst_2.INIT_RAM_31 = 256'hFC0FFCE3F98FE9113C1CFFD7FB99F0193FE7FCFBFFFFFFFFFF8FFFFF3F7FFFFC;
defparam prom_inst_2.INIT_RAM_32 = 256'hF8FF80FFFFFFFFFFF3FFFF5FD3FFFFA2477FFFFFFFFFFFFFBE3FAB5FF0BFFCE5;
defparam prom_inst_2.INIT_RAM_33 = 256'h23FFFFFFFFFFFFAFCFEBCFE67FF3837F86BF857EEFF8ADCE6B5FFBFD6EBC804F;
defparam prom_inst_2.INIT_RAM_34 = 256'hDF8D6FD7FDF7E9D737FC7F968F4E3FFD27DEBFFFFFFFFFF8FFFFF3FDFFFFFFAC;
defparam prom_inst_2.INIT_RAM_35 = 256'hE867FFFFFFFFFF9FFFF87FFFFFFF77FF0FFFFFFFFFFFE3CBF242F7977E1B9F4F;
defparam prom_inst_2.INIT_RAM_36 = 256'hFFFFFFFFFFFDFE7D983CEF3FF6A7DF9FFE87F2BFBFD87C33FF2FEF0FDC47FFC1;
defparam prom_inst_2.INIT_RAM_37 = 256'h13FDDFECF4189F7FCFFC70FF0BFFEC760DFFFFFFFFFFF3FFFFFF8FFFFEC80009;
defparam prom_inst_2.INIT_RAM_38 = 256'h7FFFFFFFFFFBFFFFFEE2FFFFF000035FFFFFFFFFFFFF3FA9EF9F8FF3FEF99FF9;
defparam prom_inst_2.INIT_RAM_39 = 256'hFFFFFFFF9FF5CB4BCEF5FC13FF7F3FB0BF1BF9FE06EEBFF9FFCA1CBDFFF51DF8;
defparam prom_inst_2.INIT_RAM_3A = 256'hA2FE1FD7D217F17F2B17416F013F8607FFFFFFFFFFBFFFF219FFFFFBFFFF313F;
defparam prom_inst_2.INIT_RAM_3B = 256'hFFFFFFFF07FFFEC797FFFE800013BFFFFFFFFFF7FBB4DBF37B7E8D3CE7DFC1EF;
defparam prom_inst_2.INIT_RAM_3C = 256'hFFFFFDFEACDE3C6EFFE7730B8BE62FE61FFA83FD67FFCFD0C9E451C835C015FF;
defparam prom_inst_2.INIT_RAM_3D = 256'hFD17FD9C3FEFFC9378747CFA75FCFFFFFFFFFFF3FFFF8BD8FFFFFFFFFFF9FFFF;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFFFCFFFFD0FFFFFFFBFFFF1BFFFFFFFFFF7E7B97EF41E7FF6BCFE3FF69FF7F;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFDFD0E0EBE109FF21B45BBE46FFA7FE449EDE0FD5FDD75E4E1DC61E8D1FFFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b1;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hC79297F1FF78030DF33FDFFF1FFFFFFFFFFF8FFFF43D4FFFFD3FFFFCBFFFFFFF;
defparam prom_inst_3.INIT_RAM_01 = 256'hFFB9FFFFDE47FFFFEBFFFEECFFFFFFFFFFF7FCCEF8907E2BBDF6DFC75FF0FFCF;
defparam prom_inst_3.INIT_RAM_02 = 256'hF97D437E345FB09F3BD5FFF3FF5FF460FE25FE3FE593F53FD7B7EF6DFFFFFFFF;
defparam prom_inst_3.INIT_RAM_03 = 256'hEFFFFFFFE3FFFFFBFFFFFFFFFFFFFFFFF57FFFF3D3FFFFE87FFFFBFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_04 = 256'h3FFFF1FFBFFFF81FFFFC57FFFFFFFE3FFFBC7FFEFFFF3FCFFFFFFFFFFFFF14FF;
defparam prom_inst_3.INIT_RAM_05 = 256'hFFFFFF0FFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFFE3F6FFFFE87FFFF37FFFFFFFFEFFF;
defparam prom_inst_3.INIT_RAM_07 = 256'hFFFFE3FFFFC3FFFFD1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFF;
defparam prom_inst_3.INIT_RAM_09 = 256'hFEE0DFCEF79F6FFCFFFFFFFFFFFBDFFFF3FE7FFFF47FFFEDFFFFFFFFFDFFFFFF;
defparam prom_inst_3.INIT_RAM_0A = 256'hFE7FFFFCBFFFFBBFFFFFFFFFFFFFB39EF7FFFFFFFFFFFC6E1FFFECEFFE00FFE4;
defparam prom_inst_3.INIT_RAM_0B = 256'hF3EFFFBFFFAF5B87BFF90D7E0033F13EB834601967CBFF3FFFFFFFFFFFA7FFFB;
defparam prom_inst_3.INIT_RAM_0C = 256'hFF633E1B93FBE7FFFFFFFFFFEFFFFC5F47FFFFCFFFFFF7FFFFFFFFEFFBA8E698;
defparam prom_inst_3.INIT_RAM_0D = 256'hFFFFE5FFFFFCFFFFFFFFFBFED61D47BD6DFF3CDDE3D6FB9FFC879F9FFFFCBF9E;
defparam prom_inst_3.INIT_RAM_0E = 256'h7FEC3738F5BFBFFF4027E00380E10B0FE1C58FEA7F65FFFFFFFFFFFEFFFFE7EE;
defparam prom_inst_3.INIT_RAM_0F = 256'h3B937D8E7CFFFFFFFFFFFFAFFFD4FBFFFFFBFFFFFF5FFFFFFFFFFFB2C726F9FF;
defparam prom_inst_3.INIT_RAM_10 = 256'hFEBFFFFF47FFFFFFFF3FE0E812593FBFFCD8315C0EFDFFF581FFFEBFA7C4CCF1;
defparam prom_inst_3.INIT_RAM_11 = 256'hE673B623A37BFB2F7FF7C9F833FCB8A6385FEB9FFFFFFFFFFFFFEFFFF6DED7FF;
defparam prom_inst_3.INIT_RAM_12 = 256'hA3CFEF4FFFFFFFFFFFFA7FFDA7B7FFFF8FFFFFC3FFFFFFFFDFF0966820E3D7FF;
defparam prom_inst_3.INIT_RAM_13 = 256'hFFFFF47FFFFFFFE7FDF52378466DFFBBE689E1F3F9FF7F5FF6B17FE70F3C5B1C;
defparam prom_inst_3.INIT_RAM_14 = 256'h20E5FD1CBE24D7EB01DFBBE31B027D2BF97907FFFFFFFFFFFD7FFFF1FF7FFFE3;
defparam prom_inst_3.INIT_RAM_15 = 256'h7739FFFFFFFFFFFF1FFFFC7FFFFFFBFFFFFFDFFFFFFFFDFF7510DE897DAFE63F;
defparam prom_inst_3.INIT_RAM_16 = 256'hFFD7FFFFFFFF3FFF7A6FABD76BF46DB0BCCF302F897DF8EB10CFCCC9CB36805E;
defparam prom_inst_3.INIT_RAM_17 = 256'h9DF92FFAEB3F49078BC2BC8DCBB24373A13FFFFFFFFFFFEAFFFFCFFBFFFEBFFF;
defparam prom_inst_3.INIT_RAM_18 = 256'h2EFFFFFFFFFFF33FFFC3FFFFFFAFFFFFF1FFFFFFFFBFFEF0938F0BDBFD2FBB2E;
defparam prom_inst_3.INIT_RAM_19 = 256'hFFFFFFFFDFFE14EEEE9BF03FDD15E79769F3FEFAFFDFE01935EFADE434DCD535;
defparam prom_inst_3.INIT_RAM_1A = 256'hA0FFC687EDDC161E1FB19B1E65F358597FFFFFFFFFFDEFFFFEBF9FFFF7FFFFF8;
defparam prom_inst_3.INIT_RAM_1B = 256'hFFFFFFFFFFE3FFFF5FEDFFF9FFFFFF9FFFFFFFC2FF9601FB898E8FC40FD7E98D;
defparam prom_inst_3.INIT_RAM_1C = 256'hFFFFF7BFFE08DF2E435FEB020DBA0E917FE897FF1FC61FFEE386EB95FCBE8E4F;
defparam prom_inst_3.INIT_RAM_1D = 256'hFCAB7FE5F7C3E37081326C0759D313FFFFFFFFFFFCFFFFCFF17FFF9FFFFF1FFF;
defparam prom_inst_3.INIT_RAM_1E = 256'hFFFFFFFFBFFFF8FD5FFF67FFFFF5FFFFFFFD1FFF7A7D9E74D0FC2827BE0AE03F;
defparam prom_inst_3.INIT_RAM_1F = 256'hFE97FFFE1EE3837E9FC3DBDFDEE65BFF0F1FF05D16FCFE80FE3E43ED5789FFFF;
defparam prom_inst_3.INIT_RAM_20 = 256'h97FF8F13FEEABB15AEC67F027D7FFFFFFFFFFFF7FFFF3EF7FFC1FFFFABFFFFFF;
defparam prom_inst_3.INIT_RAM_21 = 256'h7FF00EFFFFFFA7FFEDFFFFFCBFFFFFFEA7FFE7FFBD908FA8B893E2E39991BFF7;
defparam prom_inst_3.INIT_RAM_22 = 256'hFFFDABD225F7E6A6EC6C3EEC82FFF6E5FFF3E84FA24B15052399B7E37FFFFFFF;
defparam prom_inst_3.INIT_RAM_23 = 256'hFFF7FBE4E72E0B8F6F42CFFFFFFFFFCABC01BFFFFEFFFFB8FFFFF84FFFFFFF8B;
defparam prom_inst_3.INIT_RAM_24 = 256'hF12BFFFECB00063FFFFE55FFFFFFC7FFFF8B7288F5BE7BF8380EF57E23FEF97F;
defparam prom_inst_3.INIT_RAM_25 = 256'h0A39975C69E757FAE3C959A8FF49CFFF1E02BF3A3259E5B3F883EBFFFFFFF801;
defparam prom_inst_3.INIT_RAM_26 = 256'h7C8FAF70FEAC05F5F0FBFFFFFFFCE80021FFFFAE7FFF5FFFFFF1FFFFFFFC3FFF;
defparam prom_inst_3.INIT_RAM_27 = 256'h7FFFEDFFFF97FFFFE6FFFFFFFFAFFFE5FB6D9C1B18CBA67CF2E7CD3FFC97FF86;
defparam prom_inst_3.INIT_RAM_28 = 256'hED0702CEAA09EEDDC4D0BFFC23FFF687F3EAF97D7B633EFCBC4FFFFFFFBBFFF6;
defparam prom_inst_3.INIT_RAM_29 = 256'hFCAFB6AE4ADE9E9FB3FFFFFFDD00024FFFFDE0007BFFFFF7FFFFFFDF9FFFFDA5;
defparam prom_inst_3.INIT_RAM_2A = 256'hFFEFFFFFFFFFF99FFFFFFE1FFFFFD4BD960132FC584FBF1C00EBFF667FFEE640;
defparam prom_inst_3.INIT_RAM_2B = 256'hDE1E7A1F6763D7A399FF973FFE91C23CC0394437B15F6FF0FFFFFFFFFFFFFBFF;
defparam prom_inst_3.INIT_RAM_2C = 256'h7F786EBBDFDAEABFFFFFFFFFFFFFFFFFCFFFFFFFFFF63FFFFFFEA8FFFFD37F24;
defparam prom_inst_3.INIT_RAM_2D = 256'h7FFF80000279FFFFFF753FFFE98FC65823FED7D35E67DCBAFFE90FFFDC1FFE02;
defparam prom_inst_3.INIT_RAM_2E = 256'hE9B0E85E1CF28BEFF8F1FFEF5FFFE21F87133B1477B14FFFFFFFFFFFFFFFFFF2;
defparam prom_inst_3.INIT_RAM_2F = 256'hFCFBF13F1C67FFFFFFFFFFFFA7FFFFFFFFDFFFFF3E7FFFFF691FFFF87BFF6A07;
defparam prom_inst_3.INIT_RAM_30 = 256'hF807FF93FFFFF8EBFFFFFF5E7D38FF738AF0479FFF29F7FEFFFFF81FFCF18FEA;
defparam prom_inst_3.INIT_RAM_31 = 256'hFEE7FFFF37FFFFDFFFFFFFFFFFFFFDFFFFFEFFFFBFFFFFFFFFFFFFF7FFFFCFFF;
defparam prom_inst_3.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFBFFFF1000001E00FFFFFF8E6FFFFFFFFFFBFFFFFFF;
defparam prom_inst_3.INIT_RAM_33 = 256'h87FC7DFC0186BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE7FFFFFFE83B;
defparam prom_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFF9FFFFFE1060E6180E090100847FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_36 = 256'h0003CA1741FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFF980FFFFF0;
defparam prom_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFF1BFFFE0FFFFFFBFFFE0100FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCBFFFE5FFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3B = 256'hFFFFFFFFFFFFFC7FFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEFFFE5FFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFE7FFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b1;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7F3BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_01 = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FF;
defparam prom_inst_4.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFD883FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF97FD33F;
defparam prom_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF3FFC27FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFF;
defparam prom_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFCFFFC1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFD7FFFFFF;
defparam prom_inst_4.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFBFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFE7FFEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFF4FFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFFFEBFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFF3FFFDFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFF77FFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE2FFFFEFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1B = 256'hFFFFABFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1E = 256'hFEFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFF2FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_21 = 256'hFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;
defparam prom_inst_4.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_24 = 256'hFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF;
defparam prom_inst_4.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFE7;
defparam prom_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF7FFFF97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFF7FFF;
defparam prom_inst_4.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFF7FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFF7FFFFFFFF;
defparam prom_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFA7FFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFCFFFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFDFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5FFFFFBFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3B = 256'hFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFDFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3E = 256'hFFFF3FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b1;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE9FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_01 = 256'hE7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_04 = 256'hFFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDF;
defparam prom_inst_5.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_07 = 256'hFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFF;
defparam prom_inst_5.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFE7FFF;
defparam prom_inst_5.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFF8FFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFEFFFFFFF;
defparam prom_inst_5.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF7FFFFFFFFF;
defparam prom_inst_5.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_18 = 256'hFFFFFFFFFFFE7FFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1B = 256'hFFFFFFFFF9FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFCFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1E = 256'hFFFFFFDFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFEBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_21 = 256'hFFFDFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_24 = 256'hC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5FFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_27 = 256'hFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF;
defparam prom_inst_5.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2A = 256'hF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFF;
defparam prom_inst_5.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF83FFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2D = 256'hFFFFFE1FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF9F;
defparam prom_inst_5.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFF9D0FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_30 = 256'hFF96481A3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFDFFFFF7FFFF;
defparam prom_inst_5.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFEFFFFFE7FFFFF97FFE90FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_33 = 256'h000398FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9C000000000007FFFFFF800039C;
defparam prom_inst_5.INIT_RAM_35 = 256'h7FFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC32BFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_36 = 256'hFFF627FFFFF7E4FF7CBFFFFFF43FBFE5FFFFBFFE77B9DE7DDFC3F1FFFE7EC3FB;
defparam prom_inst_5.INIT_RAM_37 = 256'hFFCFC3361D58DE5DF07027FDAFFEDFD7FFA8000000000000FFFFFFFFFE3FFFFF;
defparam prom_inst_5.INIT_RAM_38 = 256'hB9FFFFFFFFFFFFDFFFFF90006FFFFFFFFEA8BFFFFEFB5FFC0F7FF5FFF7FFFBBF;
defparam prom_inst_5.INIT_RAM_39 = 256'hFF1FFFFF1FB3BE0FEFFD7C9CF8FF7BFBE1F38A098BBA21FCF823FAA61F97D3FF;
defparam prom_inst_5.INIT_RAM_3A = 256'hEC834060CE885A0D17BFF8D7DE7FFFFC8000000000000BFFFFE3FFFB7FFFFFFF;
defparam prom_inst_5.INIT_RAM_3B = 256'hFFFFFFFFFFFCFFFFFE0003AFFFFFFFFFA0FFFFC7F3E9C139FF5F77BEFF24FE7B;
defparam prom_inst_5.INIT_RAM_3C = 256'h3EFFFBE7BF813EFFB7E0BF57B93FCE9F6DE0AA7C7FCCE89B8DE3FEF76F8FFF87;
defparam prom_inst_5.INIT_RAM_3D = 256'h2C2848800327F06FF9BEBBFFDBFFF0000000000000BFFFFFFFFF497FFFFFFFFB;
defparam prom_inst_5.INIT_RAM_3E = 256'hFFFFFFFFD7FFFFDFFFFD7FFFFFFFFFF7FFFDBCAFEC17FFF3F97FD9FB1FFFDFE2;
defparam prom_inst_5.INIT_RAM_3F = 256'hFF3EA2FBF2C7FE5F79F0FF6DF97FFF5FF6F6E377C7DFE1FEE5BE9CF7FFFFFFFF;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b1;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h3FBF7DF9F2FA6F9ED763E7FFFFFFFFFFFFFFFFF9FFFFF3FFFFB7FFFFFFFF9D7F;
defparam prom_inst_6.INIT_RAM_01 = 256'hFFFFFEFFFFFCFFFFE9FFFFFFFFFF6FFFEFDEFEFF11FFF7CF9E7F1EFEFC3FDFFE;
defparam prom_inst_6.INIT_RAM_02 = 256'hE137BF9E3FC8F7FF9FCF9FDFFFFDFF9F5F5F3E3B7F90EF5248879FFFF3FFFFFF;
defparam prom_inst_6.INIT_RAM_03 = 256'hC3CFA7FDD7BDF6DBF5E5FFFC0000000000BFFFFFFE1FFFFFDFFFFFFFFFE3FFFE;
defparam prom_inst_6.INIT_RAM_04 = 256'h9FE7FFFFF7FFFF8FFFFFFFFFFABFFE7FD1EC7D6FF174D1EF7FFFFBFBFF3EF1E7;
defparam prom_inst_6.INIT_RAM_05 = 256'hE319C3FCFF4D7913FDFF78FF7FBC717ED6EABA77C23F9E7B78FFFF53FFF7FFFC;
defparam prom_inst_6.INIT_RAM_06 = 256'hDE3A82A29EF5897F7FFFF7FFFDFFFFFDFB7FFFFCFFFFFFFFFFFFFFFF4FFFBF37;
defparam prom_inst_6.INIT_RAM_07 = 256'h2BFFFF7FFFFFFFFFFFFFFFE1FFF3C28CD9AEFED9864E53C07F7FBFF3F9FFDEBD;
defparam prom_inst_6.INIT_RAM_08 = 256'h02BFDCF7B7DDFF1FEFDFF8FC36EFFFC7EB708DF7EB1D77CFFFF0FFFE3FFFFC7F;
defparam prom_inst_6.INIT_RAM_09 = 256'h2FEF55FFA11DF3FFFF000047FFFF5FC7FFFFDFFFFFDFFFFFFFFFF7BFFAF2AE3C;
defparam prom_inst_6.INIT_RAM_0A = 256'hFFFBFFFFF9FFFFFFFFFDBFFF5DB42D75A7E53F7EFBB94FF9FBFF3FC8FDF9CBE5;
defparam prom_inst_6.INIT_RAM_0B = 256'h8EB3DFFB03BEFF3C7F9EFD78BF79BAD2F8EB7BB3453D3FFFDFFFEFFFFFE7FEFF;
defparam prom_inst_6.INIT_RAM_0C = 256'h5D7FD65B371FFFF80003BFFFFCFEFFFFFEFFFFFCFFFFFFFFFF7BFFCF8F1BFF27;
defparam prom_inst_6.INIT_RAM_0D = 256'h8FFFFFBFFFFFFFFFFC7FFDFFF8FFACEE7EFFDFD2DFFF8F8FE9FF0F4FFF6EB8FF;
defparam prom_inst_6.INIT_RAM_0E = 256'hD5E12273D7EFCFFC7FE6E3FFF89F5FAFDFF59D25FFFFFFFFFFE7FFFF7FD7FFFF;
defparam prom_inst_6.INIT_RAM_0F = 256'hEB9F4EF8FFFFFFFFFFFFFFFFFBFFFFF37FFFE5FFFFFFFFFFFFFC7BFBBFE15BD1;
defparam prom_inst_6.INIT_RAM_10 = 256'hFFFBFFFFFFFFFFF3FF4FBDCFFDF6B7B5F8576B7DFC79FFDFF8B3FDFCBBF5EFE1;
defparam prom_inst_6.INIT_RAM_11 = 256'h13E908FF087FF7DFBC9E6380F789FD7F79D7B8FFFFFFFFFF7FFFFCFFFFFFFCDF;
defparam prom_inst_6.INIT_RAM_12 = 256'h7EE6BFFFFFFFFFEFFFFFBFBFFFFFF7FFFF3FFFFFFFFFFCFFED7FBBC1F54C796F;
defparam prom_inst_6.INIT_RAM_13 = 256'hEFFFFFFFFFFF8FFC3D76F79E061FFBE4FF465FD2DFF7F5FFCFBFF7BB3E5D3F3E;
defparam prom_inst_6.INIT_RAM_14 = 256'h21DFF393FEBE07FFF64BD7FE3FDBC72EBF3BFFFFFFFFF9FFFFCFEBFFFFF7FFFF;
defparam prom_inst_6.INIT_RAM_15 = 256'h90FFFFFFFFFEBFFFF1F5FFFFF9FFFFF3FFFFFFFFFFE5FE11FD3E9BE0D7BC7DDF;
defparam prom_inst_6.INIT_RAM_16 = 256'hFFFFFFFFFF7FF32FCFA17765FEDEFFEA2BFFA9FFEFCCFDFDBE7DC3F3FFF4DFAD;
defparam prom_inst_6.INIT_RAM_17 = 256'hFF877FEFC7BF1CF06476977E7EBEF3AA3FFFFFFFFFDFFFFAFDBFFFFF7FFFFCFF;
defparam prom_inst_6.INIT_RAM_18 = 256'hFFFFFFFFFBFFFF9F7FFFFF9FFFFFBFFFFFFFFFFF2FFB3FFFD7BE1CFDFFD1F9B4;
defparam prom_inst_6.INIT_RAM_19 = 256'hFFFFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1A = 256'hE7FFDFFFEBFFFFFFFDF3FFFDFFFFFFFFFFFFFFFDFFFFEFC5FFFFF7FFFFCFFFFF;
defparam prom_inst_6.INIT_RAM_1B = 256'hFFFFFFBFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1C = 256'hFFFEBFFFFFFFFCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFBFAFFFFFDFFFFEFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1E = 256'hFFFDFFFFDFE3FFFFEBFFFFBFFFFFFFFFFFDFFFFFFFFFD3FFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1F = 256'hFDFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFF7FCFFFFFDFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_21 = 256'hE7FFFFEF3FFFFEFFFFE7FFFFFFFFFFFE7FFFFFFFDCFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_22 = 256'hFFFFFFFF1FFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFDFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_23 = 256'h4FEC07DBD7D827FEBF903FFFFFFFFFFBFFFFBBF7FFFFEFFFF9FFFFFFFFFFFFDF;
defparam prom_inst_6.INIT_RAM_24 = 256'hFFE6F8FFFFFFFFFE5FFFFFFFFFFFFAFFF9F0FF61FFE53FC75FF01FE1CFECFFFC;
defparam prom_inst_6.INIT_RAM_25 = 256'hAF7FC077D3AFF5FBFBF3FF85FD8FFDECFDFDF9E3F5F5FF8FFFEFFFFFFFFFFF7F;
defparam prom_inst_6.INIT_RAM_26 = 256'hF87C9A7E017FF9F801FFFFFFFFFFAFFFFFFF7FFFFEBFFE5FFFFFFFFFFFFEFDB9;
defparam prom_inst_6.INIT_RAM_27 = 256'hBFDFFFFFCFFFDFFFFFFFFFFFFFDF9F67FFE2C7F7F3FAEF7E04F843FF31FFA0FC;
defparam prom_inst_6.INIT_RAM_28 = 256'hF80DFDF9FE39BF7F1FEB7F499FA70FCFEE4F9F5EBBF9BD7B7FFFFFFFFFF3FFFF;
defparam prom_inst_6.INIT_RAM_29 = 256'h8AFFF7C7FEDF8F9FFFFFFFFFFCFFFFFFFBFFFFCBFFD3FFFFFFFFFFFFDFCFFDCB;
defparam prom_inst_6.INIT_RAM_2A = 256'h7FFFF67FFDFFFFFFFFFFFFF9F1FD4B7F60FFDB1FD64FDF47D56FCDAFE473C633;
defparam prom_inst_6.INIT_RAM_2B = 256'hEFDFE5EFE9F59FEFA7FC1FF9C7FAB4FB8FF021FFAFEF5BFFFFFFFFFF3FFFFAFC;
defparam prom_inst_6.INIT_RAM_2C = 256'hBE857FF1FE20FFFFFFFFFFFFFFFEFF1FFFFFDFFDFFFFFFFFFFFFFE7FBF669FDE;
defparam prom_inst_6.INIT_RAM_2D = 256'hFFC3F27FFFFFFFFFFFFFEF4FEDDFEDDFF7FF7DF4FC1178C7FE213F493F463E5E;
defparam prom_inst_6.INIT_RAM_2E = 256'hF7FE99DFE11FD3FFBF1FCB0FFFFFEF6FC1AFFC7F80BFFFFFFFFFFFFFFF97EFFF;
defparam prom_inst_6.INIT_RAM_2F = 256'hFBFF2FFF1FFFFFFFFFFEBFFFF7FDFFFFF4FD3FFFFFFFFFFFFFF7C7FC25FFFB7E;
defparam prom_inst_6.INIT_RAM_30 = 256'hDF3FFFFFFFFFFFFFFDF1FFAEFF9C1FB39FD72FEEDFF2FFCED3F4F7FFFFFFDFD7;
defparam prom_inst_6.INIT_RAM_31 = 256'hF06BFBFFFEDFEFFBF9D6FFEFFF3DFCE1FFEBFDD3FFFFFFFFFFDFFFFE7EDFFFFF;
defparam prom_inst_6.INIT_RAM_32 = 256'hF5FF47FFFFFFFFFFEBFFFFEFF7FFFFF10F7FFFFFFFFFFFFF3E1FF7BFBFC7E66F;
defparam prom_inst_6.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFBFFCF7FFC1FC48FEFAFE7E7F6BF8DF3EEEBFF3FEEE7F3ABF;
defparam prom_inst_6.INIT_RAM_34 = 256'hFFEEFFF6FE5FEFB80FF97FF20FFEBFFE1FBEBFFFFFFFFFFD7FFFE7F4FFFFF1D3;
defparam prom_inst_6.INIT_RAM_35 = 256'hF8AFFFFFFFFFFF3FFFFAFEBFFFFE7000FFFFFFFFFFFFFBCDFFC9FFFC7EA0BFA7;
defparam prom_inst_6.INIT_RAM_36 = 256'hFFFFFFFFFFFCFF7E953F5EBF809FF213E0F3F93FE7E7FCC5FEDFF14BF013FFC7;
defparam prom_inst_6.INIT_RAM_37 = 256'hF1FEDFE5F9FD587FF7FF65FFF5FFF1FFE1FFFFFFFFFFE7FFFF3FEFFFFFE80007;
defparam prom_inst_6.INIT_RAM_38 = 256'h7FFFFFFFFFFAFFFFCFFFFFFFF7FFF87FFFFFFFFFFF7FFF660F2B9FF8B9FFE3FA;
defparam prom_inst_6.INIT_RAM_39 = 256'hFFFFFFFFFFEFFDEBE9EFFC947DB83FFE3FA7FD7C3FCE7FF1FF0A3FFE7FF9FFFC;
defparam prom_inst_6.INIT_RAM_3A = 256'hC1FFA7B7D9FFFD3FECD7BF0FFE9F7C7FFFFFFFFFFF3FFFFFFD3FFFFD0000D7FF;
defparam prom_inst_6.INIT_RAM_3B = 256'hFFFFFFFF9FFFFE3FF7FFFF00004D7FFFFFFFFFFFFBFFFEFC327E6FDFBF8FFF2F;
defparam prom_inst_6.INIT_RAM_3C = 256'hFFFFFFF9FE1C3FCA5FEFD7C39FF04BFD7FC225FB67FECFE7C1F01DF82FE84FFF;
defparam prom_inst_6.INIT_RAM_3D = 256'hFC73FC3AFFDFF776FFF274EFFDE57FFFFFFFFFF1FFFF8FD1FFFFEFFFFD3BFFFF;
defparam prom_inst_6.INIT_RAM_3E = 256'hFFFFFF7FFFE3F0FFFFF9FFFFFFFFFFFFFFFFFF0F335FF257F17AF67CF872FE27;
defparam prom_inst_6.INIT_RAM_3F = 256'hFFFFF3D0FFFDEDFA5EFDB85E44FFEFFE1F7FC76FFBFEBD1F017F80FE007FFFFF;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b1;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h7FFBEFFCFFB79FEDBFEFDFFFFFFFFFFFFFFF1FFFFF7F2FFFFFBFFFFB3FFFFFFF;
defparam prom_inst_7.INIT_RAM_01 = 256'hFFC3FFFFFF8FFFFFFFFFFF54FFFFFFFFF7E9F3FEFEB3FF1CFFDF47FFCFF0FFC9;
defparam prom_inst_7.INIT_RAM_02 = 256'hFF7E7FBFF37FDF67EDF3FFF7FF3FF2FFFF64FF5FE7FFFD3FEBA7F767FFFFFFFF;
defparam prom_inst_7.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFCBFBFFFFE3FFFFF5FFFFFFFFFD;
defparam prom_inst_7.INIT_RAM_04 = 256'h3FFFF9FEFFFFFEFFFFFD77FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF87FF;
defparam prom_inst_7.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF8FFFFF5FFFFFDFFFFFFFFFEFFF;
defparam prom_inst_7.INIT_RAM_07 = 256'hFFB7E3FFFFC7FFFFF9FFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF;
defparam prom_inst_7.INIT_RAM_09 = 256'hFDFFFFFFFFFFFFFFFFFFFFFFFFFD3FFFFDF8FFFFF9FFFFFCFFFFFFFFFDFFFFFF;
defparam prom_inst_7.INIT_RAM_0A = 256'hFF9FFFFFDFFFFFDFFFFFFFFF7FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_0B = 256'hFFFFFFFFFFFFBFFFFFFFFBFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFF8FFFF9;
defparam prom_inst_7.INIT_RAM_0C = 256'hFF9FFFFFFDFFFFFFFFFFFFFFF3FFFCFFC7FFFFF7FFFFF7FFFFFFFFEFFFDFFFFF;
defparam prom_inst_7.INIT_RAM_0D = 256'hFFFFEFFFFFFDFFFFFFFFF3FFEBFFBA7EFFFFFFFFFFEFFFFFFFFBFFFFFFFFFFFD;
defparam prom_inst_7.INIT_RAM_0E = 256'hFFF3FFC7F9FF0FFFDF1FF7FABE6E0FC37FD6FDF4FAFFFFFFFFFFFFFDFFFFFBFA;
defparam prom_inst_7.INIT_RAM_0F = 256'hCF6DFCFF1BFFFFFFFFFFFFBFFFF1FE3FFFFFFFFFFFFFFFFFFFFFFFBF38F9863C;
defparam prom_inst_7.INIT_RAM_10 = 256'hFFFFFFFFEFFFFFFFFE7FFFF6ADB01FDFFB3FCEBE7FDBFFFEF7F9FF9FFFBFFDE6;
defparam prom_inst_7.INIT_RAM_11 = 256'h3FCC0F17EB5FF8EDFF9A6E16E33F7873AF1FEF803FFFFFFFFFFFE7FFFF1FDFFF;
defparam prom_inst_7.INIT_RAM_12 = 256'h3BD6EFCFFFFFFFFFFFFBFFFFFFFBFFFFDFFFFFFDFFFFFFFFFFF1F0C7E9F9CFFC;
defparam prom_inst_7.INIT_RAM_13 = 256'hFFFFFCFFFFFFFFEFFD9FFEFA38FDFF7BDF87B3F4C2FFDF3F859D88BE4F9C5D65;
defparam prom_inst_7.INIT_RAM_14 = 256'hF1EF7C7EFFE62FECFBBEB143E3CE5CABF479F3FFFFFFFFFFFE3FFFFBFD7FFFF7;
defparam prom_inst_7.INIT_RAM_15 = 256'hCFC2FFFFFFFFFFFFF7FFFFBFFFFFFDFFFFFF1FFFFFFFFBFFDF3836F71EBFCAFB;
defparam prom_inst_7.INIT_RAM_16 = 256'hFFF7FFFFFFFFFFEDE26DFA273FF3DFA9BD0F9EBFF5A7FD104F39F0FBF4F3523C;
defparam prom_inst_7.INIT_RAM_17 = 256'h67D47FFBF9FF7FDFDF59FCF3BAEEBFA981BFFFFFFFFFFFF5FFFF2FEFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_18 = 256'h17FFFFFFFFFFFE7FFFFFFFFFFFCFFFFFFFFFFFFFFF5FFDF0FF28E9E3FFBF2E8F;
defparam prom_inst_7.INIT_RAM_19 = 256'hFFFFFFFFCFFFFE994B84B8FF66C3FFDF7D57FEFD3FFCFEFC7DFFBFCC39DFEAF9;
defparam prom_inst_7.INIT_RAM_1A = 256'hE9FFE757FFBFACBFFBF5D77F1DFCDF87BFFFFFFFFFFFBFFFFFFFBFFFF7FFFFFF;
defparam prom_inst_7.INIT_RAM_1B = 256'hFFFFFFFFFFF7FFFF9FD5FFFBFFFFFF7FFFFFFFFBFFAD4E90E9BEBFD9FE2AF3FB;
defparam prom_inst_7.INIT_RAM_1C = 256'hFFFFFBFFFFE1767C4F27FAEE257F9FE33FE6E5FFE7F30797FBFACFD43BE3637F;
defparam prom_inst_7.INIT_RAM_1D = 256'hFD797FDF7F71FDFF9D72F01E844A7FFFFFFFFFFFFEFFFFFFFD7FFE7FFFFFD7FF;
defparam prom_inst_7.INIT_RAM_1E = 256'hFFFFFFFF3FFFF8FF5FFFFFFFFFF7FFFFFFFF2FFD6DE55E72FDFB318FFFBFEE6F;
defparam prom_inst_7.INIT_RAM_1F = 256'hFF9BFF5BFAF3C12C7FDF6FDFF65FEDFF2B3FFC7EA0797F9F7DBFC5C37D87FFFF;
defparam prom_inst_7.INIT_RAM_20 = 256'hCFFFCFF29EAFE08B8750E2DF7AFFFFFFFFFFFFCFFFFF7F57FFF7FFFFFCFFFFFF;
defparam prom_inst_7.INIT_RAM_21 = 256'hFFFFF7FFFFDFAFFFF9FFFFEB3FFFFFFFCFFFDAA740E00AD9FD5DA6E266987FC2;
defparam prom_inst_7.INIT_RAM_22 = 256'hFFFEF5CFFE1ECDAEDFFD1FF7EDEFFDFFFFFBF7A783BCBD6FD49ABB813FFFFFFF;
defparam prom_inst_7.INIT_RAM_23 = 256'hFAFFFCF1FF2E38F6EE9F3FBFFFFFFFF37FFEFFFFF60FFFFE7FFFFF3FFFFFFFF3;
defparam prom_inst_7.INIT_RAM_24 = 256'h0057FFFF7B001E7FFFFF9DFFFFFFFFFFFE3B395FF563D99DE2CF906EABFE7C3F;
defparam prom_inst_7.INIT_RAM_25 = 256'hA85E369F9E53403BE1FC7E89FFD04FFF7F7E7E7BC3E15D4D800FFFFFFFFFFF2E;
defparam prom_inst_7.INIT_RAM_26 = 256'hE23FCE8AE2F64AADF7F7FFFFFFFF44005FFFFF807FFFEFFFFFFBFFFFFFFAFFFF;
defparam prom_inst_7.INIT_RAM_27 = 256'hFFFFF800007FFFFFFBFFFFFFFFBFFFDC5B87EFAF2B82157FFE3793FFEDBBFFC3;
defparam prom_inst_7.INIT_RAM_28 = 256'hFD3D1DEF795F0FBA75F97FFF28FFE4E8C7F3C6FE3533B8FDFDFFFFFFFF440008;
defparam prom_inst_7.INIT_RAM_29 = 256'hF8E7BE0A5BE31E0FAFFFFFFFF300063FFFFCE00069FFFFF9FFFFFFFEAFFFF8E6;
defparam prom_inst_7.INIT_RAM_2A = 256'hFFDFFFFFFFFFEF5FFFFFFFDFFFFF6E7E2F393E0DF063FB5F7E53FF5AFFF93FD1;
defparam prom_inst_7.INIT_RAM_2B = 256'hE1EC034FDBE2CFFF22FFEA7FFFDF3FBDFDFFCFB1F4978BF7FFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_2C = 256'h7FD73ECD77E3F1FFFFFFFFFFFFFCFFFFFFFFFFFFFFFC67FFFFFF81FFFFE81F03;
defparam prom_inst_7.INIT_RAM_2D = 256'h000060000599FFFFFF82FFFFF637FBA7DF4EF3DBB979F55ABFF0B7FF87DFCF0C;
defparam prom_inst_7.INIT_RAM_2E = 256'hF36FF43F5E7BFD7FFFFFFFFAF003C7E07FFFCFC97E7EBFFFFFFFFFFFFE7FFFF2;
defparam prom_inst_7.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003000006F7FFFFFAAFFFFFF43F9FDFD;
defparam prom_inst_7.INIT_RAM_30 = 256'hFDFFFFFFFFFFFF207FFFFFFFFEFFFFFFFFFF9FFFFCDFFFFF7FFFFFFFFFFFFFF7;
defparam prom_inst_7.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFF;
defparam prom_inst_7.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFC197FFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_33 = 256'h87FC7DFC010BDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFBFF83B;
defparam prom_inst_7.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFE3FFFFFE060E6180000FEFE07FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_36 = 256'hFFF835E93FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF63FFFFFEF;
defparam prom_inst_7.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFF3BFFFF0FC00007FFFE0101FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDEFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3B = 256'hFFFFFFFFFFFFFBBFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3E = 256'hFFFFFFFFFF8FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b1;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDF8BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_01 = 256'hDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF97DE;
defparam prom_inst_8.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE7D81FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FF8FF;
defparam prom_inst_8.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFDFFD8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFF;
defparam prom_inst_8.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFF8FFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFF9FFFFFFF;
defparam prom_inst_8.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFDFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBBFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFD7FFECBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_12 = 256'hFFFFFFFFFFFFE3FFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFE3FFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_15 = 256'hFFFFFFFFFFBFFFDCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF7DFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_18 = 256'hFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1B = 256'hFFFFABFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFBFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1E = 256'hFEFFFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFE7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_21 = 256'hFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7;
defparam prom_inst_8.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_24 = 256'hFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFF;
defparam prom_inst_8.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFF3;
defparam prom_inst_8.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFEFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF3FFF;
defparam prom_inst_8.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFEFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFDFFFFFF;
defparam prom_inst_8.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFE7FFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFCFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFBFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFA7FFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_35 = 256'hFFFFFFFFFFFF9FFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFEBFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_38 = 256'hFFFFFFFFFDFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3B = 256'hFFFFFFEFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFD3FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3E = 256'hFFFEFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b1;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFE9FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_01 = 256'hF3FFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_04 = 256'hFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F;
defparam prom_inst_9.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_07 = 256'hF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFF;
defparam prom_inst_9.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFEF;
defparam prom_inst_9.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFEFFFF;
defparam prom_inst_9.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFF;
defparam prom_inst_9.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFEFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFF7FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_18 = 256'hFFFFFFFFFFFF3FFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1B = 256'hFFFFFFFFF1FFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1E = 256'hFFFFFF9FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_21 = 256'hFFFEFFFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF3FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_24 = 256'hCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_27 = 256'hFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2A = 256'hF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFF;
defparam prom_inst_9.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFDBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2D = 256'hFFFFFFE01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFBF;
defparam prom_inst_9.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFD7FFFFD7FFFFFFD1E5FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_30 = 256'h01E479732FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0000000000005FFFFFE0000;
defparam prom_inst_9.INIT_RAM_32 = 256'hFFFFFFEFFFFFFFFFFFFE7FFFFEFFFFFFE7FFE46BFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_33 = 256'hFFFF980FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFBFFFFFDFFFFFFF;
defparam prom_inst_9.INIT_RAM_35 = 256'hFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC77FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_36 = 256'hFFF2F7FFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_37 = 256'hE7DFE01A0509E85FE8703FFABCF8FFDFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_38 = 256'hF80000000000003FFFFFA0005FFFFFFFFFF3FFFFFFFBDFA00EBFF3FEDFDFF93F;
defparam prom_inst_9.INIT_RAM_39 = 256'hF88FFFFFFF8FE00FDFF97F4DF6FC1FF8FBF3490F83F7807F789C3EB3DFF5FDFF;
defparam prom_inst_9.INIT_RAM_3A = 256'h7C2C41E81384191E237F8EC7C67EFFFD0000000000001FFFFFE40015FFFFFFFF;
defparam prom_inst_9.INIT_RAM_3B = 256'hFFFFFFFFFFF8FFFFFBFFFB5FFFFFFFFFE6FFFFEF95FF43F7FF9F42BEFFD3FFBC;
defparam prom_inst_9.INIT_RAM_3C = 256'hBFFFFFF03E9E887FE7F3EF6FAB1F8F1FB14F0FBA133707ADBFEFF7E34FDFFF9F;
defparam prom_inst_9.INIT_RAM_3D = 256'h181A61848731F069799CFEEBCBFFFFFFFFFFFFFFFF7FFFFEBFFF837FFFFFFFF9;
defparam prom_inst_9.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFD7FFFFFFFFFCFFFFFFFAFC81F7FF8F91BDDF66FE3CFC0;
defparam prom_inst_9.INIT_RAM_3F = 256'hFF4F41F3F4C7FD5CF8F3FCFDFDF1FF1FFEF1FD0FE3AFE67E7F8F3EFDFFFFFFFF;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b1;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'h3FFCE9F9EFFD639CFFEE7F3FFFFFFFFFFFFFFFF5FFFFFBFFFF87FFFFFFFF9C7F;
defparam prom_inst_10.INIT_RAM_01 = 256'hFFFFFFFFFFFCFFFFF5FFFFFFFFFEFFFFE7D73CFDB5FF675FBE0F7E7E1F7FE7FE;
defparam prom_inst_10.INIT_RAM_02 = 256'hFD4F3FC5BFDDFFDF93CFDFBF2FF4FFBFAF1FFF3DFF32E73ED0E78FFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_03 = 256'hC35F929E1719EFD2EFE7FFFCFFFFFFFFFF7FDFFFFE9FFFFE9FFFFFFFFFFFFFFA;
defparam prom_inst_10.INIT_RAM_04 = 256'h7FF7FFFFEFFFFFC7FFFFFFFFF97FFE7C69CE1B0FF7BBC7E47F57FDF3FFBF11D3;
defparam prom_inst_10.INIT_RAM_05 = 256'h6B47F7FD0EE6FAFFFBFE78FF8FC7F8F3FDECEF89A7FB9F6FFBFFFF8000000000;
defparam prom_inst_10.INIT_RAM_06 = 256'hFE0DE2FCCEA98B3F1FFFE7FFFFFFFFEFFC7FFFFBFFFFFEFFFFFFFFFFC7FFFF99;
defparam prom_inst_10.INIT_RAM_07 = 256'hDBFFFFFFFFFE7FFFFFFFFFE1FFF1C34AC8BAFF6BCE5EC7EA7FCFBFE3E0DEDFFE;
defparam prom_inst_10.INIT_RAM_08 = 256'h1E3FAC774BB6F4BFFFFFFFFA67FF8FDFFE387C23EF61CFC7FFF9FFFFFFFFFC7F;
defparam prom_inst_10.INIT_RAM_09 = 256'hCDEFD0E7C19FF1FFFE00007FFFFFDFF7FFFFCFFFFFCFFFFFFFFFF73FFE71D6B4;
defparam prom_inst_10.INIT_RAM_0A = 256'hFFFDFFFFFDFFFFFFFFFDE7FF5F3C0EF987FFCDFEE5DB3FF4E7FFFEE3EDE3EFEB;
defparam prom_inst_10.INIT_RAM_0B = 256'hDDB71FFFD79F7FFCFF8FFDFCF97EB9EBFCFE3FCF6FBEFFFFE00013FFFFF3FAFF;
defparam prom_inst_10.INIT_RAM_0C = 256'h3F0EFAFFBF0FFFFFFFFCFFFFFEFF7FFFFC7FFFFFFFFFFFFFFF73FFDFEFD3FFBB;
defparam prom_inst_10.INIT_RAM_0D = 256'hFFFFFFDFFFFFFFFFFFBFF7FBDAFF8EF365FF8F02C75FDFBFFFFF2F0E5FFF3C7E;
defparam prom_inst_10.INIT_RAM_0E = 256'hD9F7A3FDDFE9E3FF7FEFD7DFED9E5FD7A3965EE3E7FFFFFFFF97FFFF7FC7FFFF;
defparam prom_inst_10.INIT_RAM_0F = 256'hFD8F1D7DFFFFFFFFFFFFFFF7FDFFFFE3FFFFFDFFFFFFFFFFAFFEF972BFE75998;
defparam prom_inst_10.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFDFFCE1E6FFC47E63C3A6833F9F878FFBFFEFFF1FDE7EFFFE0;
defparam prom_inst_10.INIT_RAM_11 = 256'h7DE8867F143FCFFFDF7CBF1AEFB9F9BCEDF2543FFFFFFFFFFFFFFDFE7FFFFEFF;
defparam prom_inst_10.INIT_RAM_12 = 256'h7BFDEFFFFFFFFFCFFFFF3FFFFFFFFFFFFFBFFFFFFFFFFEFFFE97B3FFD3B9F8DE;
defparam prom_inst_10.INIT_RAM_13 = 256'hCFFFFFFFFFFFAFFCCFFCF7C6A27FB3C77C765FCFEFFEF22787CB087EFC3FAFDD;
defparam prom_inst_10.INIT_RAM_14 = 256'hAAEFF0B7FF3FE5FBCB3D4FC9BFC7F3BF353FFFFFFFFFF1FFFFCFFFFFFFF7FFFF;
defparam prom_inst_10.INIT_RAM_15 = 256'hB5FFFFFFFFFF3FFFF3FDFFFFFFFFFFFFFFFFFFFFFFFFFFA27DBF7BD38FAAFB3F;
defparam prom_inst_10.INIT_RAM_16 = 256'hFFFFFFFFFF7FFEFF8F207BE3F27FD7EE79FEB5FF9F2DFFFFBE67E271FDFACBDF;
defparam prom_inst_10.INIT_RAM_17 = 256'h7FF87FE3D03F3F6813FDA07F7FFDE7EDFFFFFFFFFFAFFFFE7FFFFFFE7FFFFFFF;
defparam prom_inst_10.INIT_RAM_18 = 256'hFFFFFFFFFBFFFFBFEFFFFFCFFFFF7FFFFFFFFFFFBFFFFFE7C07FCAF8AFBFFCCA;
defparam prom_inst_10.INIT_RAM_19 = 256'hFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFE7FBFFFFF3FFFFEFFFFF;
defparam prom_inst_10.INIT_RAM_1B = 256'hFFFFFF9FFFFCFF7FFFFFFFFFF3FFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1C = 256'hFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF3F8FFFFFDFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1E = 256'hFFFCFFFFFFFFFFFFE7FFFE7FFFFFFFFFFFE7FFFFFFFFA7FFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1F = 256'hFBFFFFFFFFD3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFF7FCFFFFFAFFFFDFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_21 = 256'hFFFFFF7FBFFFFE3FFFE7FFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_22 = 256'hFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_23 = 256'h47EC0FDF8FE82FFF1FD01FFFFFFFFFFBFFFFAFE7FFFFF7FFF3FFFFFFFFFFFF8F;
defparam prom_inst_10.INIT_RAM_24 = 256'hFFEFF9FFFFFBFFFC5FFFFFFFFFFFFFF5FD79FFA7FF5E3F8FDFD01FA1DFFFFFF8;
defparam prom_inst_10.INIT_RAM_25 = 256'h1DFFE37FCF1FFDC7F00FE80BF85FFE03F403E8F9FC05FFDFE01FFFFFFFFFFE7F;
defparam prom_inst_10.INIT_RAM_26 = 256'h7FB879FCFFFFFFFFFBFFFFFFFFFF9FFFFFFF3FFFFFFFFF7FFFFFFFFFFFFDFC7F;
defparam prom_inst_10.INIT_RAM_27 = 256'hBFCFFFFF8FFFCFFFFFFFFFFFFF3F2FF96FEBBFFEFBFAFFFFFDF9FEFC8CFFFF7F;
defparam prom_inst_10.INIT_RAM_28 = 256'hFEF9FF7DFFDD5F40FF97BFBEFFF8BF981FDA7F213FF9FE857FFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_29 = 256'hEE47D7EFFE8F8FFFFFFFFFFFF9FFFFDFFFFFFFD3FFC3FFFFFFFFFFFFCFE7FE77;
defparam prom_inst_10.INIT_RAM_2A = 256'hFFFFF6FFF9FFFFFFFFFFFFFDF5F8FD7E797FAFDFDF37EFFFFE3FC48FEE43EABF;
defparam prom_inst_10.INIT_RAM_2B = 256'hDFC3F7F5FDFE71FA9BF969FA32F521F9E1FBC3FFE3F897FFFFFFFFFFBFFFFDFD;
defparam prom_inst_10.INIT_RAM_2C = 256'hFEF0FFFAFFFFFFFFFFFFFFFFFFFEBFDFFFFF3FF5FFFFFFFFFFFFFE7DFFAF9FC1;
defparam prom_inst_10.INIT_RAM_2D = 256'hFFF7FA7FFFFFFFFFFFFF9F8FF6EFE603FD99F877FCFE79FEFC15FEDA3FFBFFAD;
defparam prom_inst_10.INIT_RAM_2E = 256'hEB7FE6BFBEFFDFFFBEAFDF1FFA7FEAEFFF9FFCBFFEFFFFFFFFFFF7FFFF8FE7FF;
defparam prom_inst_10.INIT_RAM_2F = 256'h7FFF8FF08FFFFFFFFFFFFFFFF1FBFFFFF9FD7FFFFFFFFFFFFFF7CFFFCBFF60FD;
defparam prom_inst_10.INIT_RAM_30 = 256'h9F3FFFFFFFFFFFFFFCFBFFF37E3EBFB9DFE9E7F9F7FA7F8797FBF3FE5FF8DFF4;
defparam prom_inst_10.INIT_RAM_31 = 256'hE40BFBDFFFFFF3F6F8237FFFFF91FDE5FFE7FDE3FFFFFFFFFFDFFFFFFF7FFFFF;
defparam prom_inst_10.INIT_RAM_32 = 256'hF4FF45FFFFFFFFFFF7FFFF9FEFFFFFC91F7FFFFFFFFFFFFFFD9FFD7FAFEFFE4F;
defparam prom_inst_10.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFCFA7FCF7FFE7FAFFFEFB7F7FFF9FF87CBF53FFE5FFC77F3B3F;
defparam prom_inst_10.INIT_RAM_34 = 256'hAFA0BFFBFEBFC7FCA7FEFFFFDFE1DFFD3FE07FFFFFFFFFFCFFFFEFF1FFFFFDD7;
defparam prom_inst_10.INIT_RAM_35 = 256'hE00FFFFFFFFFFF5FFFFFFEFFFFFF8FFFFFFFFFFFFFFFF7F1FE89FFF8FF637FD9;
defparam prom_inst_10.INIT_RAM_36 = 256'hFFFFFFFFFFFDFC7FFA7F5E1F880FD003FCB7FEFF9BE9F493FEFFFD5BFC3FFF27;
defparam prom_inst_10.INIT_RAM_37 = 256'h04FE6FF4FA7F98FFDBFFE3FE02FFC9FC33FFFFFFFFFFDFFFFF5F9FFFFFF7FFFF;
defparam prom_inst_10.INIT_RAM_38 = 256'h7FFFFFFFFFF9FFFFF7EFFFFFFFFFFCFFFFFFFFFFFF7E3FF27FF797E63FF505FE;
defparam prom_inst_10.INIT_RAM_39 = 256'hFFFFFFFFDFCFFC9FF4DFFD1FFFFDFFF9BFD3FB5FDF6E5FF7FFD8FFFDFFFEFFFE;
defparam prom_inst_10.INIT_RAM_3A = 256'hE4FF5F7FF9A7F93FD52FFFFFFEFFFF9FFFFFFFFFFF7FFFFBFCFFFFFC00015FFF;
defparam prom_inst_10.INIT_RAM_3B = 256'hFFFFFFFFFFFFFF3F77FFFF400053FFFFFFFFFFF7E1FF3DFFBE7EEC3FAF6FFE7F;
defparam prom_inst_10.INIT_RAM_3C = 256'hFFFFFDFDFFEFBFD3FF9D9FC1B7E073F97FC057FA69FF9FFECFF82FF877E07FFF;
defparam prom_inst_10.INIT_RAM_3D = 256'hF8FBFCFDFFFFFB9F7F0A7F0FFC0FFFFFFFFFFFFFFFFFCFF9FFFFF7FFFE3BFFFF;
defparam prom_inst_10.INIT_RAM_3E = 256'hFFFFFEFFFFF3FDFFFFFFFFFFBBFFFFFFFFFF7F7FF32FDE57F5CDF5ECFF87FF2F;
defparam prom_inst_10.INIT_RAM_3F = 256'hFFDFEFF4EFF763FFFC7E5FBE7BFFF9FF527FAF1FF3FF765F3E9FBB7FFA7FFFFF;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b1;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'hBFDFD3FCBFD7A7FDB7DFFFBFBFFFFFFFFFFFDFFFFE7F2FFFFEFFFFFF3FFFFFFF;
defparam prom_inst_11.INIT_RAM_01 = 256'hFFEFFFFF9FCFFFFF9FFFFF7CFFFFFFFFF7FEF934FF91FE1C5FE7DFFFCFF07FEB;
defparam prom_inst_11.INIT_RAM_02 = 256'hFEBEBEBFD6BFE7DFE1CBE803FDFFF937F0F9FFDFF2EBFEC1FC57E88FFFFFFFFF;
defparam prom_inst_11.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFBFFFFF3FFFFFBFFFFFFFFFD;
defparam prom_inst_11.INIT_RAM_04 = 256'h7FFFF9FCFFFFFDFFFFFF77FFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FCFFFFFFFFFFFAFFFFFFFFFCFFF;
defparam prom_inst_11.INIT_RAM_07 = 256'hFFFFF7FFFFF7FFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FF;
defparam prom_inst_11.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFBFEFFFFF9FFFFFD7FFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_0A = 256'h7F5FFFFFFFFFFFDFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFB;
defparam prom_inst_11.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF3FFFCFFF7FFFFBFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_0D = 256'hFFFFF3FFFFFAFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_0E = 256'hFFFFFFFFFFFF2FFF8F3FF80700F007E7EEFEFFFAFBFBFFFFFFFFFFFF7FFFEBF8;
defparam prom_inst_11.INIT_RAM_0F = 256'hFE3E7EFE81FFFFFFFFFFFFFFFFF5FF3FFFFFFFFFFFBFFFFFFFFCFFDFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_10 = 256'hFF3FFFFFCFFFFFFFFE3FEFCF7E6FEF3FFCFFF1FF7FC7FFFBFFFC00F05C3FFCDF;
defparam prom_inst_11.INIT_RAM_11 = 256'h0FD01F4FF65FFA7BFE6F83EA7DFDB3F9968FB7E0FFFFFFFFFFFFE7FFFF3FEFFF;
defparam prom_inst_11.INIT_RAM_12 = 256'hA3F5F06FFFFFFFFFFFFCFFFFF7F3FFFFDFFFFFF3FFFFFFFF9FFCF8DE9E01E3FD;
defparam prom_inst_11.INIT_RAM_13 = 256'hFFFFFCFFFFFFFFE7FFFC2DEF0371FF87F63FFDFAD7FE38BFA69F09E57FECBCFA;
defparam prom_inst_11.INIT_RAM_14 = 256'h71FEFC13FFA7BFFD407DA5DFE7F660DAF2FCDFFFFFFFFFFFFF7FFFFBFE7FFFF7;
defparam prom_inst_11.INIT_RAM_15 = 256'h5FCD7FFFFFFFFFFFC7FFFF3F9FFFFDFFFFFFDFFFFFFFFFFF8F4FBA903EBFEEFC;
defparam prom_inst_11.INIT_RAM_16 = 256'hFFEFFFFFFFFEFFF7E66E21BFEFFB9E41FA4F3ABFF1F7FE8BC00F2FF55B9F0B7F;
defparam prom_inst_11.INIT_RAM_17 = 256'h63D4EFFAF3FF84701A9C7FFB7DC3BF43FFDFFFFFFFFFFFF7FFFFBFEFFFFF3FFF;
defparam prom_inst_11.INIT_RAM_18 = 256'hDFFFFFFFFFFFFE7FFFF7FFFFFFFFFFFFF9FFFFFFFF9FFE77DBDE19E7FDBF00AE;
defparam prom_inst_11.INIT_RAM_19 = 256'hFFFFFFFFEFFF5EFD77FA77FF3BEBCBF9F0CFFE1CDFFCFFFAFA7FB7FD7F27F1FE;
defparam prom_inst_11.INIT_RAM_1A = 256'hDBFFF7E7FF5F819EFFFDFBEF51F46ECBFFFFFFFFFFFFBFFFFEFF7FFFF7FFFFFF;
defparam prom_inst_11.INIT_RAM_1B = 256'hFFFFFFFFFFFBFFFF7FDDFFFCFFFFFFFFFFFFFFFFFFE7F59DE86EFFD93BF7E89F;
defparam prom_inst_11.INIT_RAM_1C = 256'hFFFFFBFFE5C3CD799767F72E1EFE63EABFF4F1FFC7EFFFD7FEE6E3EF5E5FF9FF;
defparam prom_inst_11.INIT_RAM_1D = 256'hFEBEFFFFFAB9F3FE1C79F8AF69ED9FFFFFFFFFFFFCFFFFEFF77FFF7FFFFFCFFF;
defparam prom_inst_11.INIT_RAM_1E = 256'hFFFFFFFF3FFFFDFDDFFFBFFFFFF3FFFFFFFF7FFE3AF25F8AFFFE87BE1E4FEF6F;
defparam prom_inst_11.INIT_RAM_1F = 256'hFF1FFFEE397BE0BEFE0FFA1FF0BB47FF9E7FFF3F817DFFF6AFDE7BACF857FFFF;
defparam prom_inst_11.INIT_RAM_20 = 256'hEFFFFFED9F9FFAFF1F6DE727F8FFFFFFFFFFFFC7FFFF7F77FFEFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_21 = 256'hFFFFFBFFFFFFCFFFF9FFFFFF3FFFFFFFE7FFE3EF1EFF5F348A3FDB74E79DFFEB;
defparam prom_inst_11.INIT_RAM_22 = 256'hFFF3EBFD3BD39EA917183D09CD1FFAFBFFE7F7B7F3FF3EE1C61B3CBFBFFFFFFF;
defparam prom_inst_11.INIT_RAM_23 = 256'hFFFFE1FCFFDDFF6A4F63BF2FFFFFFFFBBFC0FFFFFEDFFFFDFFFFFFDFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_24 = 256'hFF9FFFFEC5001EBFFFFFFDFFFFFFF9FFFD1BF44FF1F948A1DAFE3A3DC7FF1D7F;
defparam prom_inst_11.INIT_RAM_25 = 256'h3E6E9BE1DD8781BBE19C1BE4FF963FFFFF833CBC1BEEFA27B7BFD3FFFFFFFC5F;
defparam prom_inst_11.INIT_RAM_26 = 256'hDFCF4EF2C186FA3BEBF6FFFFFFFF1803D3FFFF8C7FFE0FFFFFF7FFFFFFFDFFFF;
defparam prom_inst_11.INIT_RAM_27 = 256'h7FFFF3FFFFA7FFFFEFFFFFFFFFFFFFE23FECFBA63BD177BBF7EE443FF04FFFCF;
defparam prom_inst_11.INIT_RAM_28 = 256'hFF7A1DD565C10F78F47BEFF883FFE4F83BCF83FD15AF28FA7D3FFFFFFFDBFFF7;
defparam prom_inst_11.INIT_RAM_29 = 256'hF5E00F526BC3DF9FAFFFFFFFFF00067FFFFCE0006FFFFFFC7FFFFFFF9FFFF81B;
defparam prom_inst_11.INIT_RAM_2A = 256'hFFBFFFFFFFFFF95FFFFFFFEFFFFE577F7E7E709EFD5FE63E3757FECEFFFEBC36;
defparam prom_inst_11.INIT_RAM_2B = 256'h9F9DCECF7AEB9F9CF7FFE91FFFCE80BD3E03EA7CF5D7DFDFFFFFFFFFFFFFF7FF;
defparam prom_inst_11.INIT_RAM_2C = 256'hFFFCCCBC21FBF8FFFFFFFFFFFFFFFFFFC7FFFFFFFFF887FFFFFFFFFFFFE4DF77;
defparam prom_inst_11.INIT_RAM_2D = 256'hFFFFFFFFFB1DFFFFFFEFFFFFFECFF5F81FCDA7AD7CE1EDA17FFB9FFFC3DFEFDF;
defparam prom_inst_11.INIT_RAM_2E = 256'hF87DF5BF7AFF71BFFF7FFFF1F807F3C03F178F3EFCFF3FFFFFFFFFFFFEFFFFF5;
defparam prom_inst_11.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFBFFFF7FFFE5F7FFFFF97FFFFFF47FEFDF9;
defparam prom_inst_11.INIT_RAM_30 = 256'h05FFFFDFFFFFFFDF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFE000;
defparam prom_inst_11.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFC7FFFFDFFFFFFFFFFFFFFFD51FFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_33 = 256'h87FC7DFC01DE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFBFF83B;
defparam prom_inst_11.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFE7FFFFC0060E61800000003EFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_36 = 256'hFFF80404FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF43F00001F;
defparam prom_inst_11.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFBBFFFDF00000000001FEFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEFFFFBFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3B = 256'hFFFFFFFFFFFFF1BFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b1;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1F53FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_01 = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7DE;
defparam prom_inst_12.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFD85FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFBFF;
defparam prom_inst_12.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFDFFDCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFF1FFFF;
defparam prom_inst_12.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFAFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFF8FFFFFFF;
defparam prom_inst_12.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFDFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFBBFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFEE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFBFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_12 = 256'hFFFFFFFFFFFFE3FFFE5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_15 = 256'hFFFFFFFFFF7FFFD8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF73FFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_18 = 256'hFFFFFFFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEFFFFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1B = 256'hFFFFABFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1E = 256'hFCFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFF7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_21 = 256'hFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;
defparam prom_inst_12.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_24 = 256'hFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF;
defparam prom_inst_12.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF3;
defparam prom_inst_12.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFF5FFF;
defparam prom_inst_12.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFF3FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFEFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFF3FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFB7FFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_38 = 256'hFFFFFFFFFDFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFBFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3B = 256'hFFFFFFD7FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFD3FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3E = 256'hFFFEFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b1;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEDFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_01 = 256'hFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_04 = 256'hFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDF;
defparam prom_inst_13.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_07 = 256'hFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFF;
defparam prom_inst_13.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEF;
defparam prom_inst_13.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFF9FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFAFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFF;
defparam prom_inst_13.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFE7FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFE7FFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_18 = 256'hFFFFFFFFFFFF3FFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1B = 256'hFFFFFFFFF5FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1E = 256'hFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_21 = 256'hFFF9FFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_24 = 256'hEFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_27 = 256'hFFF77FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF;
defparam prom_inst_13.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2A = 256'hF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFF;
defparam prom_inst_13.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFF;
defparam prom_inst_13.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFE1E3FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_30 = 256'h01F878F69FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000001FFFFFE0000;
defparam prom_inst_13.INIT_RAM_32 = 256'hFFFFFFE80000000000007FFFFF00000078001F93FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_33 = 256'hFFFF32F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA0000000000003FFFFFC000001F;
defparam prom_inst_13.INIT_RAM_35 = 256'hFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC4FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_36 = 256'hFFF4CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_37 = 256'hEFEFC01A0F099C5BF0E019FDDEFDE7EFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_38 = 256'hF00000000000003FFFFFDFFF97FFFFFFFFFB7FFFFFFDBFD80F7FF7FFDFE7F9FF;
defparam prom_inst_13.INIT_RAM_39 = 256'hFA5FFFFF7EFFF0F5BFFDFE7DF7FEDFFFFFFC3FF3F03EBFE7BBEBFEB33F3BFDFF;
defparam prom_inst_13.INIT_RAM_3A = 256'h7CDF82EFE9C03AEF05BFF9EFB57CFFFE00000000000017FFFFE00017FFFFFFFF;
defparam prom_inst_13.INIT_RAM_3B = 256'h000000000003FFFFFE0000EFFFFFFFFFC5FFFFC7AAFD8277FFFFA77EBF00FE3D;
defparam prom_inst_13.INIT_RAM_3C = 256'hBFFFFFE3BE40B97FD3F5EFAFD53F9F1FB7F0F31FFC1EBC807BEA7FE1AFDFFFA0;
defparam prom_inst_13.INIT_RAM_3D = 256'h7FDBB7C5FF8EBFE9F8ECFA67F7FFFFFFFFFFFFFFFFFFFFFEFFFFFB7FFFFFFFF8;
defparam prom_inst_13.INIT_RAM_3E = 256'hFFFFFFFFCFFFFFCFFFF9FFFFFFFFFF83FFFF7FBFBFDB9FFDFAE7E3F1B7E7C7FD;
defparam prom_inst_13.INIT_RAM_3F = 256'hFF7F7FEFFEEFFFBDF8FFFBE7FFFBFF9FFCFFF57FEF9FE9FE257EDEFFFFFFFFFF;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b1;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'h3F7F7DFEFFFDF78D7B873EBFFFFFFFFFFFFFFFFDFFFFFBFFFFF7FFFFFFFF9AFF;
defparam prom_inst_14.INIT_RAM_01 = 256'hFFFFFFFFFFFF7FFFF9FFFFFFFFFE7FFFEBB67BFEFFFFC7BEFD7FFFFE3C7FFFFE;
defparam prom_inst_14.INIT_RAM_02 = 256'hF5BEFFCFFFF7C7A77FDF9FEF8FFFFFFF5F187F79FF1CE33EC08FAFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_03 = 256'hC77FE8DC3778F636F3F3FFFCFFFFFFFFFE7F9FFFFEBFFFFE5FFFFFFFFFE5FFF8;
defparam prom_inst_14.INIT_RAM_04 = 256'h8FF7FFFFFFFFFFF7FFFFFFFFFA7FFE3CEFBF158FFD3EBBDFFFFFFDFBFCBE1BE3;
defparam prom_inst_14.INIT_RAM_05 = 256'h7F81E3FF9E8E77BFE3FE7CFFAFC4FCFDEBF53F8BC6BBE4BF7D7FFF7FFFFFFFFF;
defparam prom_inst_14.INIT_RAM_06 = 256'h3E39DFB9AC351F9FBFFFEFFFFFFFFFE1FD7FFFFCFFFFF8FFFFFFFFFF8FFFDF1E;
defparam prom_inst_14.INIT_RAM_07 = 256'h9BFFFFBFFFFF3FFFFFFFFFE5FFF3D7DFE7DCFFF5EE7DD7E97F5F3FE7FFFE3F7B;
defparam prom_inst_14.INIT_RAM_08 = 256'hCEFFEF78FF7DF67FD3BFFBFBFF87BF7FE4778F2BCFDCD7DFFFFBFFFFFFFFFDFF;
defparam prom_inst_14.INIT_RAM_09 = 256'h5E0FBAF351F4FBFFFFFFFF8FFFFFAFFFFFFFFFFFFFCFFFFFFFFFF73FFC79E7FB;
defparam prom_inst_14.INIT_RAM_0A = 256'hFFF7FFFFF1FFFFFFFFFDDFFFFFFFFE068FFCDD46C0FFBFFDFFFF5E11F1EFEBFC;
defparam prom_inst_14.INIT_RAM_0B = 256'hFE5FDEB6269FFFFEFFCFFC3C7AFF7BEBFFF6BBEAF7FFFFFFFFFFE9FFFFFFFCFF;
defparam prom_inst_14.INIT_RAM_0C = 256'h3DAEBDFFFF8FFFFFFFFDFFFFFEFF3FFFFD7FFFFFFFFFFFFFFF7DFFFFCFCFFE3F;
defparam prom_inst_14.INIT_RAM_0D = 256'h9FFFFFFFFFFFFFFFFE3FF5EBCFFFFFEBA4E79D81AFDF8FBFFFFFBF1F7FAEFFFF;
defparam prom_inst_14.INIT_RAM_0E = 256'hD3FF1C7BFFFBDFFE7FEBEBD7F19E7FA7FBF70EEFFBFFFFFFFFF7FFFF9FE7FFFF;
defparam prom_inst_14.INIT_RAM_0F = 256'hF38FCBFFFFFFFFFFF5FFFFF7F1FFFFE7FFFFE5FFFFFFFFFF9FFC3BF4FFFF39E6;
defparam prom_inst_14.INIT_RAM_10 = 256'hFFFCFFFFFFFFFFFBFF9FDF7FF8C7F9F678C79A77FF77FF7FF8FFFDFA6F87F7FE;
defparam prom_inst_14.INIT_RAM_11 = 256'h33FDCE7FFD7FDBE17FBEF00BF3C47BBCFAE35E7FFFFFFFFF3FFFFBFFFFFFFEFF;
defparam prom_inst_14.INIT_RAM_12 = 256'h79C1DFFFFFFFFFCFFFFFFF9FFFFFFFFFFFBFFFFFFFFFFFFFF3A7C7E150DFF6FF;
defparam prom_inst_14.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFF829FDF85FF3FEAFD4FD551FD15FFDFF97FF2CC3BF72BFAFBE;
defparam prom_inst_14.INIT_RAM_14 = 256'hD327FF7FFF3EF3E1FE7D6F7D9FEFD78EFDFFFFFFFFFFF3FFFFEFEBFFFFD7FFFF;
defparam prom_inst_14.INIT_RAM_15 = 256'h65FFFFFFFFFFBFFFFFFFFFFFFBFFFFF7FFFFFFFFFFFFFF39FD3FF58BCF9DFB9F;
defparam prom_inst_14.INIT_RAM_16 = 256'hFFFFFFFFFD7FF53F9FDEF067E27CC7F3C5FF85FFDF937E7CA1ABFE0FFAF9EF9F;
defparam prom_inst_14.INIT_RAM_17 = 256'hFFCEFFFBE05FBEB01FF980FFBE71F7DE7FFFFFFFFFBFFFFD7FFFFFFFFFFFFDFF;
defparam prom_inst_14.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFBFC7FFFFAFFFFF7FFFFFFFFFFF9FF9CFFBE01CDDFDCF55FDCF;
defparam prom_inst_14.INIT_RAM_19 = 256'hFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFEFF9FFFFF7FFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1B = 256'hFFFFFF9FFFF8FF7FFFFDFFFFF3FFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1C = 256'hFFFFFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFBFCFFFFFFFFFFDFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1E = 256'hFFF9FFFFEFF3FFFFF7FFFF3FFFFFFFFFFFC7FFFFFFFFB3FFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1F = 256'hFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FDFFFFFBFFFFDFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_21 = 256'hDFFFFEFF1FFFFE3FFFFFFFFFFFFFFFFF7FFFFFFFF93FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_22 = 256'hFFFFFFFF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_23 = 256'hBFF3FFE7FFF7DFFFFFEFFFFFFFFFFFF1FFFFDFFFFFFFEFFFFFFFFFFFFFFFFFAF;
defparam prom_inst_14.INIT_RAM_24 = 256'hFFEBFDFFFFF9FFFC5FFFFFFFFFFFF7FBFEFFFFBBFFBFFFFFBFEFFFDE3FF77FFF;
defparam prom_inst_14.INIT_RAM_25 = 256'hDFBFFAFFD7BFEFFFF7FFE7FFFEFFFEFDFFFDFFEBFFFFFFD7FFF7FFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_26 = 256'hFF7E9B7FFEFFE5FBFFFFFFFFFFFFBFFFFEFEFFFFFE7FFFFFFFFFFFFFFFFFFD7E;
defparam prom_inst_14.INIT_RAM_27 = 256'h3FDFFFFFDFFFAFFFFFFFFFFFFF7FAFB32FFBCFFEEDFC7FFDFCFDFCFCBBFE3F3D;
defparam prom_inst_14.INIT_RAM_28 = 256'hFCF3FD3BFFDDFFFFFF7FFF3EBFDFFFFFCF273FBFFFFAFEFF7FFFFFFFFFEFFFFF;
defparam prom_inst_14.INIT_RAM_29 = 256'hC2B7E8C7FFEFF09FFFFFFFFFFDFFFFDFF3FFFFD3FFF3FFFFFFFFFFFFDFC3E67F;
defparam prom_inst_14.INIT_RAM_2A = 256'h7FFFF6FFEDFFFFFFFFFFFFFFFFFD62FE66FF6FDFEFBFC06F82FFA7C7E7EFD4C3;
defparam prom_inst_14.INIT_RAM_2B = 256'h8FE6F7F5EFFC2FFAC3FCCFFE9EF862FDE3FC27FFC7F01FFFFFFFFFFF3FFFF9FF;
defparam prom_inst_14.INIT_RAM_2C = 256'h7FF07FF6FFF4FFFFFFFFFFFFFFFEFF9FFFFF1FFCFFFFFFFFFFFFFFFEBFE59FD1;
defparam prom_inst_14.INIT_RAM_2D = 256'hFFFFF87FFFFFFFFFFFFFBF5FE317FE1BF1FDFA737EF7FD7FFECF7F987EED7FC3;
defparam prom_inst_14.INIT_RAM_2E = 256'h327FDDDFC3DFFDFEFEAFE7DFFB7FEEFFE17FFC7F82FFFFFFFFFFFBFFFF9FFFFF;
defparam prom_inst_14.INIT_RAM_2F = 256'h1FFFEFE0EFFFFFFFFFFF7FFFF3FDFFFFFBFEBFFFFFFFFFFFFFF3C7FC4BF872FD;
defparam prom_inst_14.INIT_RAM_30 = 256'h23BFFFFFFFFFFFFFFEFEFFB17F3EBFBF1F97B7E0F7FFFFA7E3EBD3FE3FFC27F8;
defparam prom_inst_14.INIT_RAM_31 = 256'hFDFFFE0FFF3FE9F7FB3BFF97FF40FD06FFC3FA27FFFFFFFFFFDFFFFE7FFFFFFF;
defparam prom_inst_14.INIT_RAM_32 = 256'hF3FF47FFFFFFFFFFFBFFFFFFEFFFFFCEFF7FFFFFFFFFFFFF7DBFFE9FDF7FCB8F;
defparam prom_inst_14.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFCF37FCFFFFF3FEAFFEFBFFFFFF8FFC7EBF209FF9FFF7FFFB3F;
defparam prom_inst_14.INIT_RAM_34 = 256'hFFE1DFE3FEDF1FEB27FAFFFBCFD0AFFF3FC23FFFFFFFFFFDFFFFE3FFFFFFFDF7;
defparam prom_inst_14.INIT_RAM_35 = 256'hE03FFFFFFFFFFF5FFFFFFEFFFFFFFFFFFFFFFFFFFFFFF7F3FEADFFF87E49BFE1;
defparam prom_inst_14.INIT_RAM_36 = 256'hFFFFFFFFFFFDFB7FD2FF7FBFABBFE077ECB7FCFFE7FBF577FE9FFEE7F837FF3F;
defparam prom_inst_14.INIT_RAM_37 = 256'h17FE5FECFEFFFE7FDFFEDFFE0EFFF9F807FFFFFFFFFFE7FFFFFFBFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_38 = 256'hFFFFFFFFFFFDFFFFF7F7FFFFFC0001FFFFFFFFFFFF3E1FEC6FEFF7E7E7F514FC;
defparam prom_inst_14.INIT_RAM_39 = 256'hFFFFFFFFCFFFF8D7F6FDFF91FEF93FFFFF97FF7EBFA63FECFFB13FFE3FF97FF6;
defparam prom_inst_14.INIT_RAM_3A = 256'hF5FF576FFBD7FDBFE73FFF7FFEBFFEDFFFFFFFFFFEFFFFF9FFFFFFFCFFFE9FFF;
defparam prom_inst_14.INIT_RAM_3B = 256'hFFFFFFFFEFFFFF7F77FFFF00007BFFFFFFFFFFF3F1FDB4FEB67FE77F0ECFFFEF;
defparam prom_inst_14.INIT_RAM_3C = 256'hFFFFFCFA7FB5FF5A9F9FCFD7F7E473FF7FC0EBFEFDFF9FFA79F017F057E027FF;
defparam prom_inst_14.INIT_RAM_3D = 256'hFA60FC997FE3FDDFFE06FC19FA1FFFFFFFFFFFFBFFFFEFF1FFFFFFFFFE5BFFFF;
defparam prom_inst_14.INIT_RAM_3E = 256'hFFFFFDFFFFF3FDFFFFF9FFFFE7FFFFFFFFFF3F7F935FC4CFFDDBFF7DF805FF2F;
defparam prom_inst_14.INIT_RAM_3F = 256'hFFCF93FECFF9CFFB32FEBF3FC3BFDBFE563FF7DFFDFE4F9F80DFC3FE837FFFFF;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b1;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'hFFDD97FD3F9FB7FDB7EF9FDF9FFFFFFFFFFF9FFFFDFEAFFFFFFFFFFD3FFFFFFF;
defparam prom_inst_15.INIT_RAM_01 = 256'hFFEFFFFFFFEFFFFF8FFFFFACFFFFFFFFF3FCFDF7FFA9FFBFBFBFCFFFDFF1FFDC;
defparam prom_inst_15.INIT_RAM_02 = 256'hFEFE1D3FCFFFEB8FE7E7F80FFE3FF8FFFDF9FF2FF9E5F807F807E017FFFFFFFF;
defparam prom_inst_15.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF7F7FFFFFBFFFFF5FFFFFFFFFD;
defparam prom_inst_15.INIT_RAM_04 = 256'h3FFFF8FFFFFFFCFFFFFF77FFFFFFFF7FFFFFFFFDBFFFFFFFFFFFFFFFFFFFBFFF;
defparam prom_inst_15.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFF3FEFFFFF5FFFFFFFFFFFFFFFDFFF;
defparam prom_inst_15.INIT_RAM_07 = 256'hFFDFFBFFFFFFFFFFF5FFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFF;
defparam prom_inst_15.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFF5FDFFFFFBFFFFFDFFFFFFFFFDFFFFFF;
defparam prom_inst_15.INIT_RAM_0A = 256'h7F5FFFFE7FFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFB;
defparam prom_inst_15.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF7FFFCDFEFFFFFDFFFFFFFFFFFFFFFDFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0D = 256'hFFFFEFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_0E = 256'hFFFFFFFFFFFFA7FFFFFFFFFFFFFFFFFF9F39F3FDFC07FFFFFFFFFFFC7FFFEBFC;
defparam prom_inst_15.INIT_RAM_0F = 256'hB5BFFE7EFEFFFFFFFFFFFFDFFFF7FF3FFFFEFFFFFFFFFFFFFFFEFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_10 = 256'hFFBFFFFFDFFFFFFFFEFFF7FFFFFFFFFFFFFFFFFFFFD7FFEBFFFE01D0783DF5FB;
defparam prom_inst_15.INIT_RAM_11 = 256'hDFFF9F7FF59FFD70FF00300F00FC35E71F9FB7A0BFFFFFFFFFFFE7FFFF3FFFFF;
defparam prom_inst_15.INIT_RAM_12 = 256'hFFD9E07FFFFFFFFFFFFCFFFFE7F7FFFFFFFFFFF3FFFFFFFFBFFF7F97EFFDD7FE;
defparam prom_inst_15.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFEBDAB9E0276FF73FE37D9FE2FFE5D3FC7830C873F5CBE4C;
defparam prom_inst_15.INIT_RAM_14 = 256'h15F7FC4EFF9F1FF0C103B98FDF2E7D72F63FE3FFFFFFFFFFFF7FFFF9FCFFFFFF;
defparam prom_inst_15.INIT_RAM_15 = 256'h7FB0FFFFFFFFFFFFD7FFFFFF9FFFFFFFFFFFDFFFFFFFFDFF8F3AE4B19E3FDDF2;
defparam prom_inst_15.INIT_RAM_16 = 256'hFFE7FFFFFFFEFFF7DB993FB71FF3BDE77CFFCABFFBE3FC86603FEDF1E9F3C67E;
defparam prom_inst_15.INIT_RAM_17 = 256'h37FB0FFD75FF82380B1C7F9BF3E16FE3C05FFFFFFFFFFFFDFFFFBFFFFFFFBFFF;
defparam prom_inst_15.INIT_RAM_18 = 256'h87FFFFFFFFFFFE7FFFFFF8FFFFEFFFFFF9FFFFFFFF7FF9FDD64C0DDBFC8FB83F;
defparam prom_inst_15.INIT_RAM_19 = 256'hFFFFFFFFFFFF3C339BFAFDFF6BF7EBADF4B7FE1DBFFFBF05FD7FDEFF3A1FC1FF;
defparam prom_inst_15.INIT_RAM_1A = 256'hF9FFB7FFFFFFFDBE9FE1DF9FDEF6FF39FFFFFFFFFFFFFFFFFDFF3FFFF3FFFFFF;
defparam prom_inst_15.INIT_RAM_1B = 256'hFFFFFFFFFFEFFFFF1FFDFFFBFFFFFF3FFFFFFFF7FFAF3F84F65EBFDFFAF3E6FF;
defparam prom_inst_15.INIT_RAM_1C = 256'hFFFFF8FFFEF189BE17BFFFDFDCBF3FE23FFAE5FFEBF7A7D7FBEDE7EE7FDB877F;
defparam prom_inst_15.INIT_RAM_1D = 256'hFC3DFFF3F80DE7FE993DFC27B4F05FFFFFFFFFFFFFFFFFE7FB7FFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1E = 256'hFFFFFFFFFFFFF9FEDFFFFFFFFFF7FFFFFFFF7FFC7CF64E82FDFD1BF63FECF31F;
defparam prom_inst_15.INIT_RAM_1F = 256'hFF5FFFBF9E3FDDB8FFC377F3967947FF8EDFFE1F80FCFFC74DBD4BCDDA27FFFF;
defparam prom_inst_15.INIT_RAM_20 = 256'hBFFF8FBE1EBFE9D7D72C75BF71FFFFFFFFFFFFEFFFFFBFF7FFF7FFFFF9FFFFFF;
defparam prom_inst_15.INIT_RAM_21 = 256'hFFFFFBFFFFFFEFFFFFFFFFFEBFFFFFFFFFFFDFEF5DE8BF93DD9FC7E42E8FFFCB;
defparam prom_inst_15.INIT_RAM_22 = 256'hFFFCE1D3FC238EBD7F181E4DF4FFF9E9FFF9F83FFFFDBEFBE3DFABC33FFFFFFF;
defparam prom_inst_15.INIT_RAM_23 = 256'hFEFFE1F1FF4D9F7396C33FAFFFFFFFFFC0007FFFF1C3FFFFFFFFFF5FFFFFFFEF;
defparam prom_inst_15.INIT_RAM_24 = 256'h0FBFFFFE09001EBFFFFFDDFFFFFFF9FFFD7CFB5FFDE1CFE1C10F276EFFFC1D7F;
defparam prom_inst_15.INIT_RAM_25 = 256'hBFDF17FEFB6A4171FFBC6875FF967FFF1FFDFEFFDF6FBB6B902FCBFFFFFFFF90;
defparam prom_inst_15.INIT_RAM_26 = 256'hA1EF3E81F0D76E781DF9FFFFFFFFC003BBFFFFA28001FFFFFFEFFFFFFFFC7FFF;
defparam prom_inst_15.INIT_RAM_27 = 256'h7FFFF000007FFFFFFBFFFFFFFEFFFFE37787F83F95B07F7EF622C17FE8FFFFFF;
defparam prom_inst_15.INIT_RAM_28 = 256'hFF7AFBDBEEF35F1FF4C7DFF945FFF5E05FF382BAD3CF8FFDFC3FFFFFFFE80010;
defparam prom_inst_15.INIT_RAM_29 = 256'hF5E80F3ACDDE7EBF7FFFFFFFFB00063FFFFEE00063FFFFFF7FFFFFFFCFFFFBA7;
defparam prom_inst_15.INIT_RAM_2A = 256'hFF7FFFFFFFFFF71FFFFFFFCFFFFF537FDF02769FBEDBCE5D3947FF1A7FFE3A06;
defparam prom_inst_15.INIT_RAM_2B = 256'hA07EE63E70FDBFBFB1FFCBDFFFEFFF7EBFFFCAF6F1C7FFFBFFFFFFFFFFFFE7FF;
defparam prom_inst_15.INIT_RAM_2C = 256'h81FBBE7D75FDFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFD7FFFFFFF3FFFFDF1F87;
defparam prom_inst_15.INIT_RAM_2D = 256'h0000400002D9FFFFFFCFFFFFF9EFE7F81F9FC7EF3E67E3FDFFFE4FFFD7E03FBF;
defparam prom_inst_15.INIT_RAM_2E = 256'hF5F3FBCFBDFCFAFFFFC7FFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFF7FFFF6;
defparam prom_inst_15.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF0000080000FF7FFFFF87FFFFFF87FCFE03;
defparam prom_inst_15.INIT_RAM_30 = 256'h0600001FFFFFFFD6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFE000;
defparam prom_inst_15.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFCC1FFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_33 = 256'h87FC7DFC013F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF3FF83B;
defparam prom_inst_15.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFEFFFFFE0060E618000000000FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_36 = 256'hFFF80403FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF43FFFFFFF;
defparam prom_inst_15.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFF7BFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCEFFFFBFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3B = 256'hFFFFFFFFFFFFFDBFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3E = 256'hFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_16 (
    .DO({prom_inst_16_dout_w[30:0],prom_inst_16_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_16.READ_MODE = 1'b1;
defparam prom_inst_16.BIT_WIDTH = 1;
defparam prom_inst_16.RESET_MODE = "SYNC";
defparam prom_inst_16.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFF49FFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_01 = 256'hFFFFFFFCBFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFF81FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_04 = 256'hFFFFCBFFF9AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFE5FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_07 = 256'hFE5FFFD1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFD3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0A = 256'hFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;
defparam prom_inst_16.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF57FFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0D = 256'hFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFF;
defparam prom_inst_16.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF77FFFDF;
defparam prom_inst_16.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF5FFFF8BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9BFFFF0FFF;
defparam prom_inst_16.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFF4FFFFABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFDFFFFFF;
defparam prom_inst_16.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFE57FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD9FFFFD9FFFFFFFF;
defparam prom_inst_16.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFE27FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFBBFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1E = 256'hFFFFFFFFFFFFEFFFFF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFC7FFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_21 = 256'hFFFFFFFFFF3FFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFC3FFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_24 = 256'hFFFFFFEAFFFFDDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFF37FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_27 = 256'hFFFFFFFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFF2FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2A = 256'hFDFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4FFFFC7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2D = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3;
defparam prom_inst_16.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFABFFF77FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_30 = 256'hFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FF;
defparam prom_inst_16.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF95FFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8FFFFCF;
defparam prom_inst_16.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFA7FFFEAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFF41FFF;
defparam prom_inst_16.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFDFFFFE67FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFFF5FFFFFF;
defparam prom_inst_16.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFDFFFC77FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFCBFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFB7FFDAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_16.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_17 (
    .DO({prom_inst_17_dout_w[30:0],prom_inst_17_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_17.READ_MODE = 1'b1;
defparam prom_inst_17.BIT_WIDTH = 1;
defparam prom_inst_17.RESET_MODE = "SYNC";
defparam prom_inst_17.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_01 = 256'hFFFFFFFD7FFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFF7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_04 = 256'hFFFFFBFFFDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_07 = 256'hFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFEBFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3;
defparam prom_inst_17.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5FFF;
defparam prom_inst_17.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEF;
defparam prom_inst_17.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFBFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB9FFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFE7FFFF37FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFCDFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1E = 256'hFFFFFFFFFFFFFBFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFC7FFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFE3FFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_24 = 256'hFFFFFFF1FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3FFFFBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_27 = 256'hFFFFCFFFFD5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF37FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2A = 256'hFE7FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2D = 256'hFFFE9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7;
defparam prom_inst_17.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_30 = 256'hF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFF;
defparam prom_inst_17.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2FFFFBF;
defparam prom_inst_17.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFD7FFF;
defparam prom_inst_17.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8BFFFFFF;
defparam prom_inst_17.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFDDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEBFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFDFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_17.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_18 (
    .DO({prom_inst_18_dout_w[30:0],prom_inst_18_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_18.READ_MODE = 1'b1;
defparam prom_inst_18.BIT_WIDTH = 1;
defparam prom_inst_18.RESET_MODE = "SYNC";
defparam prom_inst_18.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFF9FFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_01 = 256'hFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_04 = 256'hFFFFFBFFFDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_07 = 256'hFE1FFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFF7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0A = 256'hFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD;
defparam prom_inst_18.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0D = 256'hFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFF;
defparam prom_inst_18.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFE7;
defparam prom_inst_18.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF5FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFF;
defparam prom_inst_18.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFBFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5FFFFCFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFCFFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFCFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1E = 256'hFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFEFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_24 = 256'hFFFFFFF3FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_27 = 256'hFFFFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE6FFFF3FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2A = 256'hFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFAFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2D = 256'hFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_18.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_30 = 256'hFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFDF;
defparam prom_inst_18.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFDFFFF;
defparam prom_inst_18.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFE7FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFEFFFFFFF;
defparam prom_inst_18.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFEFFFFDEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFBFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFBFFFECFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_18.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_19 (
    .DO({prom_inst_19_dout_w[30:0],prom_inst_19_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_19.READ_MODE = 1'b1;
defparam prom_inst_19.BIT_WIDTH = 1;
defparam prom_inst_19.RESET_MODE = "SYNC";
defparam prom_inst_19.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFEFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_01 = 256'hFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_04 = 256'hFFFFF3FFFD9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFE7FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_07 = 256'hFF1FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFEBFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0A = 256'hFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9;
defparam prom_inst_19.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0D = 256'hFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFF;
defparam prom_inst_19.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7;
defparam prom_inst_19.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF1FFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF;
defparam prom_inst_19.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFDFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFDFFFFFF;
defparam prom_inst_19.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFC7FFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1E = 256'hFFFFFFFFFFFFE7FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFDFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_21 = 256'hFFFFFFFFFF3FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_24 = 256'hFFFFFFF9FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_27 = 256'hFFFFBFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFF3FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2A = 256'hFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2D = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCF;
defparam prom_inst_19.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_30 = 256'hFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFCF;
defparam prom_inst_19.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFDFFFF;
defparam prom_inst_19.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFEFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFF;
defparam prom_inst_19.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF3FFFD9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFF7FFFECFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_19.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_20 (
    .DO({prom_inst_20_dout_w[29:0],prom_inst_20_dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_20.READ_MODE = 1'b1;
defparam prom_inst_20.BIT_WIDTH = 2;
defparam prom_inst_20.RESET_MODE = "SYNC";
defparam prom_inst_20.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDDBFFFFFFCE27FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE72BFFFFFFFE23FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFAB1BFFFFFFFFB3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFAA6FFFFFFFFFE8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFF9F2CFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_0F = 256'hFFFFFFFFFFFFE8DFFFFFFFFD5BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_12 = 256'hFFFFFFFFFFDDECFFFFFFEA3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_15 = 256'hFFFFFFFE8FFFFFFFFF8BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_18 = 256'hFFFFED0BFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1B = 256'hFFC1FFFFFFFFECFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1E = 256'h83FFFFFFFD3EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_21 = 256'hFFFFFFE7AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7F;
defparam prom_inst_20.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_24 = 256'hFFFE96BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF69FFFF;
defparam prom_inst_20.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_27 = 256'hE76BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFF;
defparam prom_inst_20.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4BFFFFFFF97;
defparam prom_inst_20.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3BFBFFFFFECFFF;
defparam prom_inst_20.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF36BFFFFFFD4FFFFFF;
defparam prom_inst_20.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF63EFFFFFEE7FFFFFFFF;
defparam prom_inst_20.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7DAFFFFFFA7FFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA5BFFFFFFB3FFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF236FFFFF9AAFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_20.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_21 (
    .DO({prom_inst_21_dout_w[29:0],prom_inst_21_dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_21.READ_MODE = 1'b1;
defparam prom_inst_21.BIT_WIDTH = 2;
defparam prom_inst_21.RESET_MODE = "SYNC";
defparam prom_inst_21.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFCFFBFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFD3FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFF7FFFFFFFFFE6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFF93CFFFFFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_0F = 256'hFFFFFFFFFFFFFC4FFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_12 = 256'hFFFFFFFFFFFDFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_15 = 256'hFFFFFFFFA3FFFFFFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_18 = 256'hFFFFFFCFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1B = 256'hFFE9FFFFFFFFD6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1E = 256'hC3FFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_21 = 256'hFFFFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD3F;
defparam prom_inst_21.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_24 = 256'hFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC4FFFF;
defparam prom_inst_21.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_27 = 256'hFD3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0FFFFFFF;
defparam prom_inst_21.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03FFFFFFFD7;
defparam prom_inst_21.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4FFFFFFFFDAFFF;
defparam prom_inst_21.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFFFFFC4FFFFFF;
defparam prom_inst_21.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEB7FFFFFFF0FFFFFFFFF;
defparam prom_inst_21.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFF3BFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCCFFFFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF33FFFFFFFBFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_21.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_22 (
    .DO({prom_inst_22_dout_w[27:0],prom_inst_22_dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_8),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_22.READ_MODE = 1'b1;
defparam prom_inst_22.BIT_WIDTH = 4;
defparam prom_inst_22.RESET_MODE = "SYNC";
defparam prom_inst_22.INIT_RAM_00 = 256'hFFFE2115CDFFFFFFFFFFE4C3EEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_06 = 256'hDE7DFFFFFFFFFFFE5EFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE6;
defparam prom_inst_22.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0C = 256'hFFFFFFFFFFA6FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC02BDEE;
defparam prom_inst_22.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_12 = 256'hFFFF370EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3695FEFFFFF;
defparam prom_inst_22.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_18 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC65D1CEFEEEFFFFFF;
defparam prom_inst_22.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFED784F84ECDEEFFE5ACFFFF;
defparam prom_inst_22.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDEFB7A252122011329FFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEFFD0ECE07F3AC5ED3FFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFEDEFFEFFCD78B8ADCA8EEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_22.INIT_RAM_36 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_23 (
    .DO({prom_inst_23_dout_w[30:0],prom_inst_23_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_23.READ_MODE = 1'b1;
defparam prom_inst_23.BIT_WIDTH = 1;
defparam prom_inst_23.RESET_MODE = "SYNC";
defparam prom_inst_23.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA09FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_01 = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD834;
defparam prom_inst_23.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF827F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC800C7F;
defparam prom_inst_23.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFA0027FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8001DFFFF;
defparam prom_inst_23.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFD00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00057FFFFFF;
defparam prom_inst_23.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFF00004FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800047FFFFFFFFF;
defparam prom_inst_23.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFE80012FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00004FFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_12 = 256'hFFFFFFFFFFFFFC00017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD00001FFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_15 = 256'hFFFFFFFFFF800025FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD800083FFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_18 = 256'hFFFFFFFE00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF100005FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1B = 256'hFFFFF40001BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1E = 256'hFF00000DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000017FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_21 = 256'h00006FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_23.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_24 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_23.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000F;
defparam prom_inst_23.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFD800000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000BFFF;
defparam prom_inst_23.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFE8000017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000003FFFFFF;
defparam prom_inst_23.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFF800000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000002FFFFFFFFF;
defparam prom_inst_23.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFF800000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000005FFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_35 = 256'hFFFFFFFFFFFF8000005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4000007FFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_38 = 256'hFFFFFFFFFD000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000BFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_3B = 256'hFFFFFFE800000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800002DFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_3E = 256'hFFFF000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_23.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_24 (
    .DO({prom_inst_24_dout_w[30:0],prom_inst_24_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_24.READ_MODE = 1'b1;
defparam prom_inst_24.BIT_WIDTH = 1;
defparam prom_inst_24.RESET_MODE = "SYNC";
defparam prom_inst_24.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000015FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_01 = 256'hF0000013FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE800003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_04 = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_24.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400002FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_07 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000;
defparam prom_inst_24.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE800003F;
defparam prom_inst_24.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000003FFFF;
defparam prom_inst_24.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFF00000DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFF;
defparam prom_inst_24.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFC000005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA00001BFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFE000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000BFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_18 = 256'hFFFFFFFFFFFF400002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000005FFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1B = 256'hFFFFFFFFF6000017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE800001FFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1E = 256'hFFFFFF800000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE800002FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_21 = 256'hFFFF000009FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_24 = 256'hC000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_27 = 256'h0008FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00;
defparam prom_inst_24.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000025FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2A = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF40000;
defparam prom_inst_24.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF400001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF700000BF;
defparam prom_inst_24.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFE000003FFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_30 = 256'hFE00780E7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFC000001FFFF;
defparam prom_inst_24.INIT_RAM_32 = 256'hFFFFFFF00000000000008000010000007FFFFD57FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_33 = 256'h000089AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFC000003FFFFFE0;
defparam prom_inst_24.INIT_RAM_35 = 256'hFFFFC000000000000000000000000000000039FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_36 = 256'h000D8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_24.INIT_RAM_37 = 256'hFFFFFFFDFEF7FFA7FFFFFFFFFFFFFFFFFFC00000000000000000000000000000;
defparam prom_inst_24.INIT_RAM_38 = 256'hF0000000000000200000400018000000001AFFFFFDFFFFFFFFFFFFFF2FFFFD7F;
defparam prom_inst_24.INIT_RAM_39 = 256'h06DFFFFFBEEFE6FBEFFFFF7BFFFD37FDF7F7FFFD7FEBFEF7FFFEFFE7FEBBF7FF;
defparam prom_inst_24.INIT_RAM_3A = 256'hFF32FD7208BFF96EFDEFDFD7FE7EFFFF00000000000010000017FFE000000000;
defparam prom_inst_24.INIT_RAM_3B = 256'h000000000001000001FFFDD00000000039FFFFCF8FFB3C63FE5FFEFEBFE9FE7F;
defparam prom_inst_24.INIT_RAM_3C = 256'hFFFFF5E7FE709FFFAFD83FCFF4FFAFDFBB20B37AE81EA1C0BBFF71E19FBFFFC0;
defparam prom_inst_24.INIT_RAM_3D = 256'h7FF7F7DC7F8FBFFCFD8F7FF7E7FFFFFFFFFFFFFFFF000001FFFFE88000000006;
defparam prom_inst_24.INIT_RAM_3E = 256'hFFFFFFFFF000000FFFFD80000000007FFFFF7DFF9FF79FEEF9F3EFE39FE7C7FF;
defparam prom_inst_24.INIT_RAM_3F = 256'hFFFEBFE7FDEFFB7C7EF87DF7FEF5FF3FF8F1F98FE3AFF3DF7F9EDEFEFFFFFFFF;

pROM prom_inst_25 (
    .DO({prom_inst_25_dout_w[30:0],prom_inst_25_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_25.READ_MODE = 1'b1;
defparam prom_inst_25.BIT_WIDTH = 1;
defparam prom_inst_25.RESET_MODE = "SYNC";
defparam prom_inst_25.INIT_RAM_00 = 256'h7D7CE7F8E3FF57DD77EEBF3FFFFFFFFFFFFFFFFE000007FFFFD80000000064FF;
defparam prom_inst_25.INIT_RAM_01 = 256'hFFFFFE000003FFFFF000000000015FFFE7FCF9FF3DFECF5EFE1FBEFFBEFFEFFE;
defparam prom_inst_25.INIT_RAM_02 = 256'hF5CE7FBDFFBBEBCF97FFBFF7DFF1FFFFDF1EFE3CFF3EF79AF7DFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_03 = 256'hEFFF977FD67DEFB479EBFFFEFFFFFFFFFEFFE000011FFFFF600000000017FFFB;
defparam prom_inst_25.INIT_RAM_04 = 256'h3FF0000007FFFFD800000000077FFE3E739FEFBFEE7F7DE3FF9FF1F3FFFFFFFF;
defparam prom_inst_25.INIT_RAM_05 = 256'hE7BD7BFBFF0079DFCFFCF8FFAFFA7AF8E7FB1FFDEFF7EECEFFFFFFC000000000;
defparam prom_inst_25.INIT_RAM_06 = 256'h7C49E3F5FEFB473F5FFFE80000000007FE800007FFFFF900000000006FFFDF7C;
defparam prom_inst_25.INIT_RAM_07 = 256'hE40000BFFFFF40000000001FFFE7F739E099FEEBDDBE67DDFF5EBFF3F0FF3F7D;
defparam prom_inst_25.INIT_RAM_08 = 256'h1EFFAD7F179DFAFFFFDFF8F817CFCFEFE1782E7FAC76FFCFFFFC00000000027F;
defparam prom_inst_25.INIT_RAM_09 = 256'hDC0BAFF3F399F9FFFE7FFFC000001FF800000FFFFFE000000000087FFCFAF278;
defparam prom_inst_25.INIT_RAM_0A = 256'h000BFFFFFE00000000023FFF1EFF9F05DFEFDFBBEEB9DFFAFDFEFF0BF3E7EDEF;
defparam prom_inst_25.INIT_RAM_0B = 256'hFAE33E3FCF7FFF7CFFD7FE7D7CFCFEE7FDF9F8FCCFBDFFFFFFFFFA000003FD00;
defparam prom_inst_25.INIT_RAM_0C = 256'hBCFFFC3B8FBFFFFFFFFF000001FFC000037FFFFF800000000089FFDFCFE7FEF1;
defparam prom_inst_25.INIT_RAM_0D = 256'h1FFFFFC000000000007FF3E3F9FFAEFEDCD79F77EF9FCF3FF7FFEFFFDF6FBBFE;
defparam prom_inst_25.INIT_RAM_0E = 256'h3BFBA0BBFFEFFFFE7FEFEFDFFB9FFFFFEFCFFD73E3FFFFFFFFE80000FFE80000;
defparam prom_inst_25.INIT_RAM_0F = 256'hFFDFDDFDFFFFFFFFFA000017FE000017FFFFFA00000000007FFF7EFC7FE79DA0;
defparam prom_inst_25.INIT_RAM_10 = 256'hFFFD00000000000DFFAF3E1FF9CE6FCF7EE79FF9FCFBFF3FFCFAF9FDF3EFF3FF;
defparam prom_inst_25.INIT_RAM_11 = 256'h59FFBD7F0FFFF7FF3E3D7F29F9FF7D7CF4E30F7FFFFFFFFE400001FF800000FF;
defparam prom_inst_25.INIT_RAM_12 = 256'hBCFF7FFFFFFFFFC000007F800000FFFFFF8000000000007FE1EF97FE7C8BF7EF;
defparam prom_inst_25.INIT_RAM_13 = 256'hC000000000004FFCEBFFF826A2FEAFE67E577FEF7FF8F81FBFFC223C619F3F7D;
defparam prom_inst_25.INIT_RAM_14 = 256'h3FC7FFDFFF3CF1FFE37BBFBDB7CFE75EBFDBFFFFFFFFFE00002FFC00003FFFFF;
defparam prom_inst_25.INIT_RAM_15 = 256'h79FFFFFFFFFF400003FF000003FFFFF8000000000003FFBDFD3DF99EAFABF7FF;
defparam prom_inst_25.INIT_RAM_16 = 256'h0000000002FFFFBF8F01773BFBFCC7EFBFFFFBFF9F417FFCC013FF83FAFBDFEF;
defparam prom_inst_25.INIT_RAM_17 = 256'hFFEEFFF7E03F7F700CFBC07E7F7BFBEEFFFFFFFFFFD00002FF800001FFFFFE00;
defparam prom_inst_25.INIT_RAM_18 = 256'hFFFFFFFFF000007FE800007FFFFF8000000000007FFDDFE7E03EDDFEDFBBFBEE;
defparam prom_inst_25.INIT_RAM_19 = 256'h00000017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000FF8000007FFFFC00000;
defparam prom_inst_25.INIT_RAM_1B = 256'hFFFFFF800005FF800002FFFFF0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_1C = 256'h0000FFFFFFFFFCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE800003FD000007FFFFF00000000;
defparam prom_inst_25.INIT_RAM_1E = 256'hFFFF00003FF000001FFFFF4000000000002FFFFFFFFF07FFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_1F = 256'h03FFFFFFFFC5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFD000005FFFFA00000000000;
defparam prom_inst_25.INIT_RAM_21 = 256'hD00000FFE000017FFFF0000000000001FFFFFFFFF83FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_22 = 256'hFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_25.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00007FE000001FFFFE0000000000007F;
defparam prom_inst_25.INIT_RAM_24 = 256'h0017F8000003FFFFA0000000000007FFFFFFFFD7FFFFFFFFFFFFFFFFFFF8FFFF;
defparam prom_inst_25.INIT_RAM_25 = 256'h3E7FE0FFEFCFF3E7F807F007FD1FFF03F803F1F7F803FFEFF00FFFFFFFFFFE00;
defparam prom_inst_25.INIT_RAM_26 = 256'h00FC3B7F007FF3FC07FFFFFFFFFFA00003FFC000007FFF40000000000003FEFF;
defparam prom_inst_25.INIT_RAM_27 = 256'hFFE000003FFFF0000000000000FF5FCB9FF78FF1C7FE70FE03FE03FF31FFC0FE;
defparam prom_inst_25.INIT_RAM_28 = 256'hFB03FC3D7FBC7F803F80BF007F800F003F461F807FFE7F017FFFFFFFFFF00000;
defparam prom_inst_25.INIT_RAM_29 = 256'hFED7FFBFFF9FFFFFFFFFFFFFFD000027F0000027FFF400000000000027D3F8D3;
defparam prom_inst_25.INIT_RAM_2A = 256'h80000AFFFA00000000000007FFFC98FE037FED5F870FEF8FD9EFC87FE3D3EF37;
defparam prom_inst_25.INIT_RAM_2B = 256'hDFCF9FFDD7F037E247E1E1FD86F843FD4FF811FFD3F027FFFFFFFFFFC00007FF;
defparam prom_inst_25.INIT_RAM_2C = 256'hFF0E7FFEFC01FFFFFFFFFFC00001FFE00000BFFF00000000000001FC7FD63FFE;
defparam prom_inst_25.INIT_RAM_2D = 256'h0017FF800000000000007F8FFA77E7B7F885FBF8FF00FE51FFB7FF64FF04FF62;
defparam prom_inst_25.INIT_RAM_2E = 256'hBFFE807FFD7FE7FF5E7FFF8FFDFFEF9FFFFFFCFFFDBFFFFFFFFFFA00004FE000;
defparam prom_inst_25.INIT_RAM_2F = 256'h67FF1FE06FFFFFFFFFFF80000FFC000007FFC000000000000007DFFF1FFAFFFC;
defparam prom_inst_25.INIT_RAM_30 = 256'h82A000000000000002F5FFD8FE7D7F5BDFC80FF0CFFD7FC7D3E7CBFE9FFDB3F8;
defparam prom_inst_25.INIT_RAM_31 = 256'hF1E5FA05FFFFF1F5FF89FFF7FFE4FE01FFF3FC1FFFFFFFFFFFA00000FF800000;
defparam prom_inst_25.INIT_RAM_32 = 256'hF7FEB8FFFFFFFFFFF400005FD0000020E080000000000000BF7FFE9FFFC7F5F7;
defparam prom_inst_25.INIT_RAM_33 = 256'h000000000000003F8FFC1FFFEBFDB3FD047F807F97FE7EFF0D7FEDFFF8FF447F;
defparam prom_inst_25.INIT_RAM_34 = 256'h3FA15FEFFEFF2FC7DFFEFFF8BFE06FFDFFC23FFFFFFFFFFD000017FA00000A18;
defparam prom_inst_25.INIT_RAM_35 = 256'hEF7FFFFFFFFFFFE00002FE00000000000000000000000FE9FFC7FFFCFE96FFF1;
defparam prom_inst_25.INIT_RAM_36 = 256'h000000000002FF7FC37FBF1FE2EFC7AFFB07F97F97C3FB19FEFFFFB3FFDFFF8F;
defparam prom_inst_25.INIT_RAM_37 = 256'hEBFFBFFBF0FC7A7F87FF33FFF1FFE3FFCBFFFFFFFFFFF00000FFE00000000000;
defparam prom_inst_25.INIT_RAM_38 = 256'hFFFFFFFFFFF800001FFC00000BFFFE800000000000BE7FFC3FC7D7E17FF9E9FF;
defparam prom_inst_25.INIT_RAM_39 = 256'h000000002F87F7EBFDEDF992FFFCFFFE7FC7FD3E3F1E7FF1FFEDFFFF3FFF7FF8;
defparam prom_inst_25.INIT_RAM_3A = 256'hFBFF7F4FC38FFEFFEB8FFF7FFEFFFF7FFFFFFFFFFF000005FD000002FFFF6000;
defparam prom_inst_25.INIT_RAM_3B = 256'hFFFFFFFFE00001FFC800003FFF9700000000000BF9FF5AFFBCFF1DFF3F1FFF3F;
defparam prom_inst_25.INIT_RAM_3C = 256'h000002FBFF6D7F471FA52FEBEBFC6FFEBFE3B7F5F5FFEFF163F82BF06FF057FF;
defparam prom_inst_25.INIT_RAM_3D = 256'hFBDCFE3AFFD3FE797C04FE11F813FFFFFFFFFFF000003FFE00001FFFFFE40000;
defparam prom_inst_25.INIT_RAM_3E = 256'hFFFFFE00000BF8000001FFFFDC0000000000BE1FCB8FFE3FEAF7F9F0F908FF4F;
defparam prom_inst_25.INIT_RAM_3F = 256'h002FC7EBFFFDF3FE38FF5EBE3C3FD7FFF5FF5EBFFFFF3FDFBF7FFDFFFCFFFFFF;

pROM prom_inst_26 (
    .DO({prom_inst_26_dout_w[30:0],prom_inst_26_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_26.READ_MODE = 1'b1;
defparam prom_inst_26.BIT_WIDTH = 1;
defparam prom_inst_26.RESET_MODE = "SYNC";
defparam prom_inst_26.INIT_RAM_00 = 256'h5FE3E7FF3FCBE7F24FF05FA03FFFFFFFFFFF800002FF5000007FFFFD40000000;
defparam prom_inst_26.INIT_RAM_01 = 256'hFFF000001FC000007FFFFF93000000000BFBFAF2FF06FFDF7F872FA00FFBFFE0;
defparam prom_inst_26.INIT_RAM_02 = 256'hFC7F3E7FE97FC7CFF3E7F007FE7FFD2FF8F3FF9FF1F3F803F00FF00FFFFFFFFF;
defparam prom_inst_26.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FF800000BFFFFFE0000000002;
defparam prom_inst_26.INIT_RAM_04 = 256'h800005FF000000FFFFFE0800000000FFFFFFFFFE7FFFFFFFFFFFFFFFFFFFCFFF;
defparam prom_inst_26.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000003F900000BFFFFF90000000002FFF;
defparam prom_inst_26.INIT_RAM_07 = 256'h000FF4000017FFFFFA000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam prom_inst_26.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE40000FFF000007FFFFFE8000000003FFFFFF;
defparam prom_inst_26.INIT_RAM_0A = 256'h7FA000007FFFFF8000000000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00005;
defparam prom_inst_26.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF400035FF800007FFFFFE8000000003FFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0D = 256'h000017FFFFFF000000000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_0E = 256'hFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800017FD;
defparam prom_inst_26.INIT_RAM_0F = 256'hCE7CFF3F01FFFFFFFFFFFFE0000BFFC00003FFFFFF0000000003FFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_10 = 256'h00FFFFFFD0000000017FFFFFFFFFFFFFFFFFFFFFFFFDFFF7CFFFFFEFBFC3FBE7;
defparam prom_inst_26.INIT_RAM_11 = 256'h1F803F1FFF3FFDFBFF00780F807DB8EBCF1F27C07FFFFFFFFFFFE000003FF000;
defparam prom_inst_26.INIT_RAM_12 = 256'hE7D5E7BFFFFFFFFFFFFF00000FF000002FFFFFF8000000007FFDFBF79A07E7FE;
defparam prom_inst_26.INIT_RAM_13 = 256'hFFFFFE000000001FFE1EE9C2FC71FFC7F9C7C3FFFFFE9EFFF87EF198DF8F3D6F;
defparam prom_inst_26.INIT_RAM_14 = 256'h6DF17EBFFFCFCFF79BFC7777DF8FB87FF5FDEBFFFFFFFFFFFF400007FE80000B;
defparam prom_inst_26.INIT_RAM_15 = 256'hFE03FFFFFFFFFFFFC80001FF800002FFFFFFA000000007FFCFCB73CEBFFFF2FB;
defparam prom_inst_26.INIT_RAM_16 = 256'hFFF8000000007FFDDBEC77D7CFFDFF46FDDF6ABFF9DBFEBFC0E9CDFAF7EF1DBF;
defparam prom_inst_26.INIT_RAM_17 = 256'h43D32FF9F7FFFCFFDBF3FE3874E46FAFFEBFFFFFFFFFFFFE00006FE00000FFFF;
defparam prom_inst_26.INIT_RAM_18 = 256'hC7FFFFFFFFFFFE000003FD00003FFFFFFE00000000FFF9FDE33FE7DBFE37875F;
defparam prom_inst_26.INIT_RAM_19 = 256'h000000003FFEDCF2CFFFFDFFCFE9FFFBF8FBFFDF7FFDBFF7FAFFF6BF3DD7E07F;
defparam prom_inst_26.INIT_RAM_1A = 256'hEBFFEFCFFFDFC17F9FE5A73FAFFCBFF3FFFFFFFFFFFF800002FF000007FFFFFE;
defparam prom_inst_26.INIT_RAM_1B = 256'hFFFFFFFFFFF40000DFE20005FFFFFF8000000007FFFF8F71FF1C7FE07EFCFD3F;
defparam prom_inst_26.INIT_RAM_1C = 256'h000007FFF1FBE478238FF0CE41B99FD9FFF5FFFFCFEFCFFFFC73F3E9BD0F877F;
defparam prom_inst_26.INIT_RAM_1D = 256'hFE3A7FF8FBF7E7FE9C77F9CF56EFFFFFFFFFFFFFFC000007F48001FFFFFFD000;
defparam prom_inst_26.INIT_RAM_1E = 256'hFFFFFFFF400005FD20001FFFFFF8000000017FFF3B6D3FFEE7FCC7DEDE73FACF;
defparam prom_inst_26.INIT_RAM_1F = 256'h00DFFFBF9CAF9FFB7F9BF1EF973983FFDEDFFFBE867B7F9F9F7EB5D67BD7FFFF;
defparam prom_inst_26.INIT_RAM_20 = 256'hEFFFB7E1DFFFF5CBAF8A71D777FFFFFFFFFFFFF800003F880017FFFFFF000000;
defparam prom_inst_26.INIT_RAM_21 = 256'hFFFFFC00003FE00003FFFFFEC00000003FFFDBBF49E0FF99EC9C7CE6DF51FFCB;
defparam prom_inst_26.INIT_RAM_22 = 256'hFFF3E3FA7FDBDFF2F779BF8397FFF6EFFFF9FFBFC7FEF0F9C9DEB7FC7FFFFFFF;
defparam prom_inst_26.INIT_RAM_23 = 256'hFBFFF7FCFF6E3F7CCFA0FFAFFFFFFFFC000100000C2C0000FFFFFFC00000001F;
defparam prom_inst_26.INIT_RAM_24 = 256'h0FA000013AFFE17FFFFFC200000001FFFFF97C3FFAE3CC0EDFB7E477DFFEF8FF;
defparam prom_inst_26.INIT_RAM_25 = 256'hD61E4FFF7C773EF3F9C39A7BFFF71FFF3FFC7EFFE787FEB5EFCFDFFFFFFFFEE0;
defparam prom_inst_26.INIT_RAM_26 = 256'hFFBF6EF0FB769D660BF3FFFFFFFFC003FC000060FFFF3FFFFFE4000000017FFF;
defparam prom_inst_26.INIT_RAM_27 = 256'h80000FFFFFDFFFFFF200000001FFFFED67DBE057D0E83CBBE41B54FFEDE7FF97;
defparam prom_inst_26.INIT_RAM_28 = 256'hFC79E7F531E9FF3AF7C29FFDBFFFF9F023CFE3FD19F7F97A7FBFFFFFFFE7FFEE;
defparam prom_inst_26.INIT_RAM_29 = 256'hFFE7EFFEE7F27FBF8FFFFFFFFB0006600003E00067FFFFFA800000007FFFFFFD;
defparam prom_inst_26.INIT_RAM_2A = 256'h00BFFFFFFFFFFBE000000067FFFF757C1E7D76FA7873969FD577FF3C7FFFFDFA;
defparam prom_inst_26.INIT_RAM_2B = 256'hFFDE9BDEDEF7E7B749FFFCBFFFDFFFBFF9FFED7A788F9FFBFFFFFFFFFFFFF800;
defparam prom_inst_26.INIT_RAM_2C = 256'h00FD5F3EFBF3FCFFFFFFFFFFFFF800003FFFFFFFFFFCF80000001FFFFFE8BFFF;
defparam prom_inst_26.INIT_RAM_2D = 256'hFFFF8000034600000031FFFFFCFFF7F017C9CFC63CF3F3D2FFFD1FFFEFE01FCF;
defparam prom_inst_26.INIT_RAM_2E = 256'hF8FFFFFFFFFFFC7FFF8FFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFF40000D;
defparam prom_inst_26.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0000080001000008080000075FFFFFF8FFFFFFF;
defparam prom_inst_26.INIT_RAM_30 = 256'h07FFFFE000000024FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF400002000;
defparam prom_inst_26.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFE8000020000000000000003CEFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_33 = 256'h78038203FEAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA00000C007C4;
defparam prom_inst_26.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFF8000020060E618000000015FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_36 = 256'h0007FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000BC0000000;
defparam prom_inst_26.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFF440002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE100003FFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3B = 256'hFFFFFFFFFFFFFC40002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE900001FFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3E = 256'hFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_26.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_27 (
    .DO({prom_inst_27_dout_w[30:0],prom_inst_27_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_27.READ_MODE = 1'b1;
defparam prom_inst_27.BIT_WIDTH = 1;
defparam prom_inst_27.RESET_MODE = "SYNC";
defparam prom_inst_27.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_01 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFF2;
defparam prom_inst_27.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFAFF;
defparam prom_inst_27.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFF7FFFF;
defparam prom_inst_27.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFDFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFF;
defparam prom_inst_27.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFDFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFF3FFFFFFFFF;
defparam prom_inst_27.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_12 = 256'hFFFFFFFFFFFFF7FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_15 = 256'hFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF3FFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_18 = 256'hFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_1B = 256'hFFFFDFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_1E = 256'hFCFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_21 = 256'hFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;
defparam prom_inst_27.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_24 = 256'hFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFF;
defparam prom_inst_27.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFBFFF;
defparam prom_inst_27.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFF;
defparam prom_inst_27.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFBFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFE7FFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_3B = 256'hFFFFFFEFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_3E = 256'hFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_27.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_28 (
    .DO({prom_inst_28_dout_w[30:0],prom_inst_28_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_28.READ_MODE = 1'b1;
defparam prom_inst_28.BIT_WIDTH = 1;
defparam prom_inst_28.RESET_MODE = "SYNC";
defparam prom_inst_28.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFDFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_01 = 256'hFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_04 = 256'hFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBF;
defparam prom_inst_28.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_07 = 256'hF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDF;
defparam prom_inst_28.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFF;
defparam prom_inst_28.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFF;
defparam prom_inst_28.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFF;
defparam prom_inst_28.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFE7FFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFDFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1B = 256'hFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1E = 256'hFFFFFF9FFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_21 = 256'hFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFF7FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_27 = 256'hFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7F;
defparam prom_inst_28.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFF;
defparam prom_inst_28.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F;
defparam prom_inst_28.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFE7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_30 = 256'h00007801FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000005FFFFFC0000;
defparam prom_inst_28.INIT_RAM_32 = 256'hFFFFFFF0000000000000FFFFFF0000007FFFFCCFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_33 = 256'hFFFF879FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_35 = 256'hFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_36 = 256'hFFFC5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_38 = 256'hFC0000000000003FFFFFC0001FFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFEFF;
defparam prom_inst_28.INIT_RAM_39 = 256'hFE7FFFFF7F77FF03DFFCFF83F9FE0FFBFBF80603807701F81C077F7FBF7DFBFF;
defparam prom_inst_28.INIT_RAM_3A = 256'hFDCFFE5CFEEFBEF7FA9FAAEF9EFD7FFE0000000000001FFFFFE00005FFFFFFFF;
defparam prom_inst_28.INIT_RAM_3B = 256'hFFFFFFFFFFFDFFFFF9FFFE9FFFFFFFFFEBFFFFEFB9FABEFBFF3F8E7D7FADFF7C;
defparam prom_inst_28.INIT_RAM_3C = 256'hFFFFFBEA3EA09DFFE7F43F0FC1BFFF3F3360BBFF7A0E65C123E2F9E79F1FFFFF;
defparam prom_inst_28.INIT_RAM_3D = 256'hFFEFDFFFFFFEFF9CFAFFFE63E7FFFFFFFFFFFFFFFFBFFFFFFFFFFBFFFFFFFFFE;
defparam prom_inst_28.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFD7FFFDFBEFAFEF7FFBF7FFD3F3EFEBF7FE;
defparam prom_inst_28.INIT_RAM_3F = 256'hFFDFF1EBFDF7FFBFF9F77EF1F8FFFF5FFFF9FFAFFFCFFF1EBB9F18FBFFFFFFFF;

pROM prom_inst_29 (
    .DO({prom_inst_29_dout_w[30:0],prom_inst_29_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_29.READ_MODE = 1'b1;
defparam prom_inst_29.BIT_WIDTH = 1;
defparam prom_inst_29.RESET_MODE = "SYNC";
defparam prom_inst_29.INIT_RAM_00 = 256'hBEFD7BFFFFFEFFACEFBFFFFFFFFFFFFFFFFFFFFBFFFFF3FFFFDFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_01 = 256'hFFFFFF7FFFFFFFFFF9FFFFFFFFFF1FFFE7EFFAFEF1FFAFFFBD3F7DFF3E7FDFFE;
defparam prom_inst_29.INIT_RAM_02 = 256'hF39EBFEEFFE5E7CF4BFF7FDF9FFFFF9FDFDDFEBCFF59EB5FE7CF8FFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_03 = 256'hFFCFFF7FC7FADF38B3F3FFFF0000000001FFFFFFFFFFFFFFFFFFFFFFFFFBFFFF;
defparam prom_inst_29.INIT_RAM_04 = 256'h5FFFFFFFE7FFFFEFFFFFFFFFFEFFFEFD73AFFFFFFB78F7D7FFCFFFE7FF7FE7EF;
defparam prom_inst_29.INIT_RAM_05 = 256'hEBC0FFFEAF5FF53FE1FD7EFF9F81FFFFFBF6D70BCE3DFD2C7DFFFF0000000000;
defparam prom_inst_29.INIT_RAM_06 = 256'h7EC9C2798E737FFFFFFFDFFFFFFFFFEBFEFFFFFFFFFFF9FFFFFFFFFFFFFF8FFC;
defparam prom_inst_29.INIT_RAM_07 = 256'hFFFFFF7FFFFFFFFFFFFFFFFFFFF3FF9AF03AFFBBF49D77EFFF9FFFEBE01F3FBC;
defparam prom_inst_29.INIT_RAM_08 = 256'h177FFDFAF759F37FEFDFFFFC27FFAFFF8EF05E639FFFF7D7FFF9FFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_09 = 256'h5FE3C8EBDBF9F5FFFF7FFFEFFFFF9FEFFFFFCFFFFFCFFFFFFFFFFE7FFCF9FEBC;
defparam prom_inst_29.INIT_RAM_0A = 256'hFFFFFFFFFBFFFFFFFFFFCFFFFE38AFFDFFFC9F03D8BEBFFFF7FFBFF7F3FFF7E4;
defparam prom_inst_29.INIT_RAM_0B = 256'hFFEFFFF1DE7FFFBE7FCFFFFFFFFC7DFFFBFE3FECD6FEFFFFFFFFF7FFFFFFFDFF;
defparam prom_inst_29.INIT_RAM_0C = 256'hFE0FBF37CFFFFFFFFFFEFFFFFCFFFFFFFEFFFFFFFFFFFFFFFFFFFFC7AF6BFEFF;
defparam prom_inst_29.INIT_RAM_0D = 256'h9FFFFF9FFFFFFFFFFE7FF9FFC2FFDF77C6FFAC818FFFAFFFF1FFDFDFBFDF7EFF;
defparam prom_inst_29.INIT_RAM_0E = 256'hF9E37FE3EFF7F7FD7FE3EFC7E3AF7FEFA3CE0FFFFFFFFFFFFFCFFFFFFFCFFFFF;
defparam prom_inst_29.INIT_RAM_0F = 256'hF1D3FDFEFFFFFFFFFBFFFFEFFBFFFFFFFFFFF7FFFFFFFFFFCFFE7EF8BFE35CEF;
defparam prom_inst_29.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFF3EEFFCFFFBD67CD7CDF9FFFBFFDFFAFDF5FC6BFFF1E4;
defparam prom_inst_29.INIT_RAM_11 = 256'hF5F7DF7F5FFFF7FEFE7FFFFFF3FC7E3FF3EF9FBFFFFFFFFFFFFFF9FFFFFFFDFF;
defparam prom_inst_29.INIT_RAM_12 = 256'hFAFB8FFFFFFFFFEFFFFFFFDFFFFFFFFFFFBFFFFFFFFFFE7FEBEFEBFF7FFEFFBF;
defparam prom_inst_29.INIT_RAM_13 = 256'hCFFFFFFFFFFFFFFF73FCFFDE3FBE7BFD7CEB9FF3BFF9FFEFEFDFE3FFFF7F2FDF;
defparam prom_inst_29.INIT_RAM_14 = 256'hDBF7FBEFFEFEFFF3EF7DFF99AFF3EF1FBBEFFFFFFFFFFFFFFFDFF7FFFFEFFFFF;
defparam prom_inst_29.INIT_RAM_15 = 256'hC7FFFFFFFFFE7FFFF3FFFFFFF9FFFFF3FFFFFFFFFFF3FF3FFEFFF7DCDFECF55F;
defparam prom_inst_29.INIT_RAM_16 = 256'hFFFFFFFFFFFFE8FF9FFFFCFFF3BE6FE747FF47FFCFFFFEF9FFB3F6FFFBFFF7CF;
defparam prom_inst_29.INIT_RAM_17 = 256'hFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFF3FFFFFFFFFFCFF;
defparam prom_inst_29.INIT_RAM_18 = 256'hFFFFFFFFF3FFFF9FFFFFFFDFFFFF3FFFFFFFFFFF9FFE3FFFFFFF3FFFFFFFFFF1;
defparam prom_inst_29.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFEFF9FFFFF3FFFFCFFFFF;
defparam prom_inst_29.INIT_RAM_1B = 256'hFFFFFF9FFFFFFE7FFFFFFFFFF3FFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFF7FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_1E = 256'hFFFFFFFFFFF3FFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFF33FFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_1F = 256'hF9FFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFBFEFFFFFFFFFFDFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_21 = 256'hEFFFFE7FFFFFFF7FFFE7FFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_22 = 256'hFFFFFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFEFFFFFFFFFFFFFFFFFDF;
defparam prom_inst_29.INIT_RAM_24 = 256'hFFF7FFFFFFFFFFFEFFFFFFFFFFFFF3FFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_25 = 256'hFFFFF1FFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7F;
defparam prom_inst_29.INIT_RAM_26 = 256'hFF7EBFFEFEFFF5FFFDFFFFFFFFFFDFFFFEFFFFFFFEFFFF7FFFFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_27 = 256'hFFCFFFFFDFFFDFFFFFFFFFFFFFBF5FDFAFF45FF5EFFAFFFDFFFBFFFECBFF7F7E;
defparam prom_inst_29.INIT_RAM_28 = 256'hFDF3FFF3FF9FBFFFFFFFFFFE7FFFFFFFFFAE1FBF9FFDFFFF7FFFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_29 = 256'hE597E027FF7FC0FFFFFFFFFFFDFFFFEFFFFFFFFFFFF7FFFFFFFFFFFFEFFFFEEF;
defparam prom_inst_29.INIT_RAM_2A = 256'hFFFFFFFFF3FFFFFFFFFFFFFDFCFF9FFE5A7FDDFF87AFD07FA31FCB4FF61FE187;
defparam prom_inst_29.INIT_RAM_2B = 256'hFFC3F7E5EFF83BF3C7FD2FFB0DFC71FDF7FC11FFFFF01FFFFFFFFFFF3FFFFDFF;
defparam prom_inst_29.INIT_RAM_2C = 256'hFFF87FFDFFFFFFFFFFFFFFFFFFFF7F9FFFFFBFF9FFFFFFFFFFFFFFFC3F9BFFB9;
defparam prom_inst_29.INIT_RAM_2D = 256'hFFEFFDFFFFFFFFFFFFFFDF0FF3EFE9F3F0FDFDFFFFFAFFFFF97F7EDC3FEFFFE5;
defparam prom_inst_29.INIT_RAM_2E = 256'hA7FF7FBFFEFFEFFE7F7FB70FFBFFF47FFE7FFC3FFF7FFFFFFFFFFBFFFFDFFFFF;
defparam prom_inst_29.INIT_RAM_2F = 256'h9FFF0FFFDFFFFFFFFFFE7FFFFBFDFFFFFDFE7FFFFFFFFFFFFFF7EFFF19FCF3FE;
defparam prom_inst_29.INIT_RAM_30 = 256'hFCFFFFFFFFFFFFFFFFFBFFF47FFFBFBB7FF06FFF3FFBFF87FFF7EBFFFFFEDFFF;
defparam prom_inst_29.INIT_RAM_31 = 256'hFC0FFFEBFEDFE1F4FF0BFFEFFFA7FFF7FFC3FFD3FFFFFFFFFFFFFFFFFF3FFFFF;
defparam prom_inst_29.INIT_RAM_32 = 256'hFBFEFCFFFFFFFFFFF7FFFFFFFFFFFFC0BFFFFFFFFFFFFFFFBEFFFE9FFFEFEFB7;
defparam prom_inst_29.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFCFFFFE9FB77FFFFFE7EFFD7F87CBFA1FFEBFFEF3FFFFF;
defparam prom_inst_29.INIT_RAM_34 = 256'hDFFEFFF7FF7FAFFFFFFA7FF2CFFF5FFEFFFC3FFFFFFFFFFEFFFFF7FBFFFFF81F;
defparam prom_inst_29.INIT_RAM_35 = 256'hF03FFFFFFFFFFFFFFFFDFF7FFFFFFFFFFFFFFFFFFFFFFBFFFF4FFFF87FC1FFEE;
defparam prom_inst_29.INIT_RAM_36 = 256'hFFFFFFFFFFFEFEFF9FFFFE1FF97FC437F03FFFFFFFEBFF1FFFDFFFD3F833FFFF;
defparam prom_inst_29.INIT_RAM_37 = 256'hFDFFDFFDFAFE87FFD7FF43FFF0FFFFFFFFFFFFFFFFFFE7FFFFBFFFFFFFFFFFFF;
defparam prom_inst_29.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFF7FFFFF80000FFFFFFFFFFFFBE1FFDDFCF97E1DBF1F5FF;
defparam prom_inst_29.INIT_RAM_39 = 256'hFFFFFFFFEF87FA77F9EDF99AFCFFFFFF7FD7FD3CBFBE1FF5FFBEFFFC3FFEFFFF;
defparam prom_inst_29.INIT_RAM_3A = 256'hF7FFAF6FEB87FDFFFDFFFFBFFE9FFFBFFFFFFFFFFF7FFFFBFEFFFFFC00005FFF;
defparam prom_inst_29.INIT_RAM_3B = 256'hFFFFFFFFCFFFFF7FFFFFFF3FFFE5FFFFFFFFFFFBE1FDFDFD7E7E66FFFFFFFF7F;
defparam prom_inst_29.INIT_RAM_3C = 256'hFFFFFEFDFFED3F52BFDBFFFFF7F47FFDFFE213FBE5FF7FFAFFF82FF027E02FFF;
defparam prom_inst_29.INIT_RAM_3D = 256'hFDAFFFFDFFFFFDFEFE07FC19FC19FFFFFFFFFFFFFFFFFFEFFFFFFFFFFF3FFFFF;
defparam prom_inst_29.INIT_RAM_3E = 256'hFFFFFEFFFFF7FFFFFFFFFFFFEFFFFFFFFFFFBFFFD70FED6FF7FBFEF5FF0FFFFF;
defparam prom_inst_29.INIT_RAM_3F = 256'hFFEFFFEFCFFBF3FD3AFFBDFFFF7FFBFF367FAF7FFCFFEFBFBFBF7FFFFE7FFFFF;

pROM prom_inst_30 (
    .DO({prom_inst_30_dout_w[30:0],prom_inst_30_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_30.READ_MODE = 1'b1;
defparam prom_inst_30.BIT_WIDTH = 1;
defparam prom_inst_30.RESET_MODE = "SYNC";
defparam prom_inst_30.INIT_RAM_00 = 256'h7FF7E7FCFFE79FE01FE01F805FFFFFFFFFFFDFFFFEFF7FFFFE7FFFFE7FFFFFFF;
defparam prom_inst_30.INIT_RAM_01 = 256'hFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFBFBF87CFF43FFAE3F9F9FE03FFCFFE0;
defparam prom_inst_30.INIT_RAM_02 = 256'hFFFFFFFFF0FFFFFFFFFFFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFE7FFFFFFF7FFFFF3FFFFFFFFFE;
defparam prom_inst_30.INIT_RAM_04 = 256'hBFFFFDFEFFFFFCFFFFFE7FFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_07 = 256'hFFCFFFFFFFEFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF;
defparam prom_inst_30.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFDFFFFF9FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_0A = 256'hFFBFFFFE7FFFFF9FFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam prom_inst_30.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFF7FFFFFFFFEFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFF9;
defparam prom_inst_30.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFCFF7FFFFDFFFFFF3FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_10 = 256'hFF7FFFFFEFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_11 = 256'hFFDFBFFFE8BFFBFDFFFFB7F6FF7FFAFDB7FF9FBFBFFFFFFFFFFFF7FFFF3FFFFF;
defparam prom_inst_30.INIT_RAM_12 = 256'hF7EDE7FFFFFFFFFFFFFDFFFFFFFBFFFFDFFFFFFFFFFFFFFFDFFBFDBF7FFFFFFE;
defparam prom_inst_30.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFEBDE9DF7EF5FFB7E7EFDBFFE7FEBDFFDFFFFD9FFF0FF96F;
defparam prom_inst_30.INIT_RAM_14 = 256'h0FF77FB5FF87FFF8C301E9CFEFAF7C77FB7A0FFFFFFFFFFFFF7FFFF9FFFFFFF7;
defparam prom_inst_30.INIT_RAM_15 = 256'hEF06FFFFFFFFFFFFEFFFFFFF9FFFFDFFFFFFFFFFFFFFFDFF87FDF7E09DFFEDFB;
defparam prom_inst_30.INIT_RAM_16 = 256'hFFFFFFFFFFFEFFE5D7DD77D7FFFBBFE77DFFB6FFE1D7FE96E0DDADFFEFDFC7FC;
defparam prom_inst_30.INIT_RAM_17 = 256'h47E3EFFFFEFFFFFFFFFBFFFFFFFD5F3FFEBFFFFFFFFFFFFBFFFFDFF7FFFF7FFF;
defparam prom_inst_30.INIT_RAM_18 = 256'h8FFFFFFFFFFFFE7FFFF3FFFFFFDFFFFFFFFFFFFFFFBFFFF4C35FFFD7FEFFAF5F;
defparam prom_inst_30.INIT_RAM_19 = 256'hFFFFFFFFFFFFFEBFD7FF74FFE9EBDFF7F9CFFFFFBFFD7FFEFAFFEFDFFCD3C0FF;
defparam prom_inst_30.INIT_RAM_1A = 256'hFAFFF7EFFF4FFFBEBFE3D70FBEF55FE1FFFFFFFFFFFFDFFFFFFF3FFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFBFCFFFFFFFFFFFFFFFFFFFF3FFF7AFB7FF5EBFFD7A7FFEBF;
defparam prom_inst_30.INIT_RAM_1C = 256'hFFFFFDFFF5EB85FBD7AFFFFFE37FD7EDFFF5EFFFEBF86F97F87FC3FDBD57BB7F;
defparam prom_inst_30.INIT_RAM_1D = 256'hFC7FFFFAFDFFFFFF1DFBFDEF5FFFFFFFFFFFFFFFFCFFFFE7FBFFFFFFFFFFEFFF;
defparam prom_inst_30.INIT_RAM_1E = 256'hFFFFFFFFBFFFFFFEFFFF9FFFFFF3FFFFFFFF7FFD7FFF7FFFEFFFE3D94FFFF7CF;
defparam prom_inst_30.INIT_RAM_1F = 256'hFFBFFF2FFC7FA1BFFF5FFFFBF57FD7FF0EBFFEBFFBFFFFFF5EFEDFD7F81FFFFF;
defparam prom_inst_30.INIT_RAM_20 = 256'hA7FFFFC1BFDFFFFFFFEBF46E7DFFFFFFFFFFFFFFFFFF7F3FFFEFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_21 = 256'hFFFFF9FFFFFFEFFFFFFFFFFF7FFFFFFFFFFFEBA78DF0BFFFDBFFC6FF6E4BFFFB;
defparam prom_inst_30.INIT_RAM_22 = 256'hFFFFF1FF7FFF85F7B7A6B96F9BFFFFFDFFFFFFF7D7FF7FFFEFBFCDFD7FFFFFFF;
defparam prom_inst_30.INIT_RAM_23 = 256'hFA7FF5F5FF5EBEF687E3FF3FFFFFFFF800017FFFF807FFFCFFFFFFDFFFFFFFF3;
defparam prom_inst_30.INIT_RAM_24 = 256'h0FBFFFFF03FFFFFFFFFFEFFFFFFFF9FFFFBD78DFFAF13D8FEFFE66E7FFFEBD7F;
defparam prom_inst_30.INIT_RAM_25 = 256'hBF5FD7FEFD437F3FFF9FDC77FFBF5FFE1FFD7CBFC3FF9FF5FFDFEBFFFFFFFF00;
defparam prom_inst_30.INIT_RAM_26 = 256'hDFFFAFF8EA2F5D7C0BFFFFFFFFFF8003FFFFFFE0FFFF5FFFFFFFFFFFFFFDFFFF;
defparam prom_inst_30.INIT_RAM_27 = 256'hFFFFF800002FFFFFFBFFFFFFFF3FFFF6F7DDF07F60F03FFA6637EBFFF677FFD7;
defparam prom_inst_30.INIT_RAM_28 = 256'hF7FE0DF73FFFEE1A7EC7DFFDEDFFF5F03FFF83FD7FBF7FFFFFFFFFFFFFF00000;
defparam prom_inst_30.INIT_RAM_29 = 256'hFEF7FF3EEDFFFE9FAFFFFFFFFCFFF9FFFFFE1FFF9FFFFFFEFFFFFFFF9FFFFFED;
defparam prom_inst_30.INIT_RAM_2A = 256'hFFBFFFFFFFFFFD7FFFFFFFCFFFFFB6FFFFFF7ACDF87BD6BEFD77FFFFFFFDFDFD;
defparam prom_inst_30.INIT_RAM_2B = 256'hE01E0F9F99F99F9E87FFE03FFF9F00FE7E07E0B9F5D7E7E7FFFFFFFFFFFFE7FF;
defparam prom_inst_30.INIT_RAM_2C = 256'hFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFE7FFFFFFFE7FFFFE03F8F;
defparam prom_inst_30.INIT_RAM_2D = 256'h00000000039FFFFFFFEBFFFFFEDFFBFFEFEBFFFFFFFFFFE1FFFE3FFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFC;
defparam prom_inst_30.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFCFFFFF7FFFE00000FFFFFFFFF7FFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_30 = 256'h07FFFFFFFFFFFFEDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_30.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFC5FFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_33 = 256'hFFFFFFFFFF99FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFDFF9F19E7FFFFFFFF3FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFF7FFFFFFFF;
defparam prom_inst_30.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3B = 256'hFFFFFFFFFFFFF9FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3E = 256'hFFFFFFFFFFDFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_31 (
    .DO({prom_inst_31_dout_w[30:0],prom_inst_31_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_31.READ_MODE = 1'b1;
defparam prom_inst_31.BIT_WIDTH = 1;
defparam prom_inst_31.RESET_MODE = "SYNC";
defparam prom_inst_31.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3F8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1;
defparam prom_inst_31.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF9FF;
defparam prom_inst_31.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFBFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFF;
defparam prom_inst_31.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFDFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFCFFFFFFF;
defparam prom_inst_31.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFF7FFFFFFFFF;
defparam prom_inst_31.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFEFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFDFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_12 = 256'hFFFFFFFFFFFFF7FFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_15 = 256'hFFFFFFFFFFBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_18 = 256'hFFFFFFFBFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_1B = 256'hFFFFDFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_1E = 256'hFEFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_21 = 256'hFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7;
defparam prom_inst_31.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_24 = 256'hFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF;
defparam prom_inst_31.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7;
defparam prom_inst_31.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_35 = 256'hFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_3B = 256'hFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_3E = 256'hFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_32 (
    .DO({prom_inst_32_dout_w[30:0],prom_inst_32_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_32.READ_MODE = 1'b1;
defparam prom_inst_32.BIT_WIDTH = 1;
defparam prom_inst_32.RESET_MODE = "SYNC";
defparam prom_inst_32.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_01 = 256'hFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_04 = 256'hFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_07 = 256'hFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFF;
defparam prom_inst_32.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDF;
defparam prom_inst_32.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFF;
defparam prom_inst_32.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFF;
defparam prom_inst_32.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFEFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFFFFF;
defparam prom_inst_32.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFF7FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_18 = 256'hFFFFFFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_1B = 256'hFFFFFFFFFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_1E = 256'hFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_21 = 256'hFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_24 = 256'hEFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F;
defparam prom_inst_32.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7F;
defparam prom_inst_32.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_30 = 256'hFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFBFFFF;
defparam prom_inst_32.INIT_RAM_32 = 256'hFFFFFFE0000000000000FFFFFF0000007FFFFC3FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_33 = 256'hFFFF807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_35 = 256'hFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_36 = 256'hFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_38 = 256'hF80000000000003FFFFFC0001FFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_39 = 256'hFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_32.INIT_RAM_3A = 256'hFE0180E01DC07C0701DFDDEFCF7EFFFFFFFFFFFFFFFFE7FFFFEFFFF9FFFFFFFF;
defparam prom_inst_32.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFBFFFF1FFFFFFFFFE7FFFFDFDDFDC0F7FF3FC0FE7F13FEFE;
defparam prom_inst_32.INIT_RAM_3C = 256'h7FFFF3F77F7F3CFFEFE39F9FCE7F9FBFC0FF1C4731FF19FE77F73BF3DFBFFFFF;
defparam prom_inst_32.INIT_RAM_3D = 256'hFFE7FFCE7F9FFFCEFDCE7AF7EFFFFFFFFFFFFFFFFFBFFFFF7FFFF3FFFFFFFFFE;
defparam prom_inst_32.INIT_RAM_3E = 256'hFFFFFFFFEFFFFFDFFFFE7FFFFFFFFFCFFFFFFCCFDFE73FF9F9E7E3F7CFF7EFFC;
defparam prom_inst_32.INIT_RAM_3F = 256'hFFFF3BF7F9CFFE7E7DF8FDFBFDF9FFBFF9FBF3DFE7DFF3BF73DE3DF9FFFFFFFF;

pROM prom_inst_33 (
    .DO({prom_inst_33_dout_w[30:0],prom_inst_33_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_33.READ_MODE = 1'b1;
defparam prom_inst_33.BIT_WIDTH = 1;
defparam prom_inst_33.RESET_MODE = "SYNC";
defparam prom_inst_33.INIT_RAM_00 = 256'h7E7EF3F9F3FCE7DEFF873E7FFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFDFF;
defparam prom_inst_33.INIT_RAM_01 = 256'hFFFFFF7FFFFEFFFFFDFFFFFFFFFF3FFFEFCE7DFFFBFFDF9FFEDFFE7F7F7FE7FF;
defparam prom_inst_33.INIT_RAM_02 = 256'hFBDF7FFE7FFBF7DFB7FF9FCFDFF9FFCF9FBE7F7EFFBDF7BFE9EFDFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_03 = 256'hE79FCFFFEF3DE77B7BF7FFFFFFFFFFFFFFFFDFFFFFBFFFFF7FFFFFFFFFF7FFF9;
defparam prom_inst_33.INIT_RAM_04 = 256'h3FFFFFFFEFFFFFEFFFFFFFFFFEFFFF7EF7DFFB9FFEFDF3ECFFE7F3F7FE7FF3FF;
defparam prom_inst_33.INIT_RAM_05 = 256'hF7FCE7FFDFBCFBBFF3FEFDFFDFFCFFF9F3F9FFF1EF79CEDEFCFFFF8000000000;
defparam prom_inst_33.INIT_RAM_06 = 256'hFF33FC7BDF7BB39F3FFFEFFFFFFFFFE7FEFFFFFDFFFFFDFFFFFFFFFFDFFFDF9E;
defparam prom_inst_33.INIT_RAM_07 = 256'hBFFFFF7FFFFF7FFFFFFFFFFBFFF7E7BDFF3DFFF7E33EEFF0FFBF3FF7FF3F7E7E;
defparam prom_inst_33.INIT_RAM_08 = 256'hFF3FFEFE1FBDFAFFE7FFFCFFCFCFDFBFC07F9F77DFCCE7EFFFFDFFFFFFFFFEFF;
defparam prom_inst_33.INIT_RAM_09 = 256'h9FF7DDF7F73DFBFFFF80000FFFFFBFFFFFFFDFFFFFEFFFFFFFFFFEFFFDFDE77F;
defparam prom_inst_33.INIT_RAM_0A = 256'hFFFBFFFFFBFFFFFFFFFFDFFF3F7DDFFFCFFB3E79E7FC7FF9FFFF3FF9FBF3F3F3;
defparam prom_inst_33.INIT_RAM_0B = 256'hFE079E780F3FFE7EFFEFFE7FFCFEF9FFFCF37CE5EFFE7FFFFFFFFBFFFFF7FDFF;
defparam prom_inst_33.INIT_RAM_0C = 256'h3EDF3979DF9FFFFFFFFF7FFFFDFF7FFFFEFFFFFEFFFFFFFFFFFBFFEFDF37FE73;
defparam prom_inst_33.INIT_RAM_0D = 256'hBFFFFFDFFFFFFFFFFEFFFBF3EDFF9CFFB9E7DE7BDFFFDF9FFBFF9FFF3F9E7FFF;
defparam prom_inst_33.INIT_RAM_0E = 256'h3DF79E77F7F3E7FEFFF7E7EFF7DF3FCF97EF5E73E7FFFFFFFFEFFFFFBFEFFFFF;
defparam prom_inst_33.INIT_RAM_0F = 256'hFBC79FF9FFFFFFFFFFFFFFEFFBFFFFF7FFFFF7FFFFFFFFFFDFFEFCFB7FF7BFFF;
defparam prom_inst_33.INIT_RAM_10 = 256'hFFFDFFFFFFFFFFFBFF9FBF1FFDE73FEF7DEFDCFDFCFFFF9FFDF9FBFEF7CFFBF1;
defparam prom_inst_33.INIT_RAM_11 = 256'h3BF33E7FBEFFE7FF3F7E7F9CFBFEFC7E71F7BE7FFFFFFFFF7FFFFBFEFFFFFDFF;
defparam prom_inst_33.INIT_RAM_12 = 256'h7DEF9FFFFFFFFFEFFFFF7FDFFFFFBFFFFF3FFFFFFFFFFEFFF7CFC7FF39CFF9FF;
defparam prom_inst_33.INIT_RAM_13 = 256'hEFFFFFFFFFFFDFFCF3F5FFCF73FF7FCEFEE79FE7BFFDFFCFFF9FF73FFF9FBF9D;
defparam prom_inst_33.INIT_RAM_14 = 256'hBC0FFC07FF7F03F7F780CFBE47E7F7BF7C07FFFFFFFFFBFFFFDFF7FFFFEFFFFF;
defparam prom_inst_33.INIT_RAM_15 = 256'h83FFFFFFFFFF7FFFF7FDFFFFFBFFFFFBFFFFFFFFFFF7FFC0FE7E03E1DFDDFBBF;
defparam prom_inst_33.INIT_RAM_16 = 256'hFFFFFFFFFEFFF07FFF80F877FF7FFFFF83FF83FFFF80FDFFC07FEF01FDFDEFFF;
defparam prom_inst_33.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEFFBFFFFF7FFFFEFF;
defparam prom_inst_33.INIT_RAM_18 = 256'hFFFFFFFFFBFFFFBFEFFFFFDFFFFFBFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_19 = 256'hFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFE7FDFFFFF7FFFFEFFFFF;
defparam prom_inst_33.INIT_RAM_1B = 256'hFFFFFFDFFFFDFF7FFFFEFFFFFBFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_1C = 256'hFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFF7FDFFFFFFFFFFDFFFFFFFF;
defparam prom_inst_33.INIT_RAM_1E = 256'hFFFDFFFFEFFBFFFFFFFFFF7FFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_1F = 256'hFBFFFFFFFFE9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFBFEFFFFFDFFFFDFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_21 = 256'hEFFFFEFFBFFFFF7FFFF7FFFFFFFFFFFF7FFFFFFFF87FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_22 = 256'hFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFDFF7FFFFFFFFFBFFFFFFFFFFFFDF;
defparam prom_inst_33.INIT_RAM_24 = 256'hFFF7FDFFFFFBFFFEFFFFFFFFFFFFF7FFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F;
defparam prom_inst_33.INIT_RAM_26 = 256'h00FF7CFF01FFFBFC03FFFFFFFFFFDFFFFFFF7FFFFEFFFFFFFFFFFFFFFFFEFFFF;
defparam prom_inst_33.INIT_RAM_27 = 256'hBFEFFFFFFFFFDFFFFFFFFFFFFFBFBFE7DFF83FFBF3FDF9FE01FC01FF07FF80FF;
defparam prom_inst_33.INIT_RAM_28 = 256'hFDF7FD7BFEBFFF7FFEFFFFBEFFDFDFBFDFAF3FFFBFFD7FFFFFFFFFFFFFF7FFFF;
defparam prom_inst_33.INIT_RAM_29 = 256'hF5DFF02FFF5FC0DFFFFFFFFFFFFFFFEFFBFFFFF7FFE7FFFFFFFFFFFFEFD7F7EB;
defparam prom_inst_33.INIT_RAM_2A = 256'hFFFFFFFFFBFFFFFFFFFFFFFFF5FEBAFF42FF5FFFCFBFE07FC31FE85FF617F18F;
defparam prom_inst_33.INIT_RAM_2B = 256'hDFE77FF7EBFFDFFCFFF4CBFF75FFEFFFB5FFE3FFD7FFD7FFFFFFFFFFBFFFFFFE;
defparam prom_inst_33.INIT_RAM_2C = 256'h7FFCFFF5FFF5FFFFFFFFFFEFFFFF7FDFFFFFFFFDFFFFFFFFFFFFFF7E7FD6BFB6;
defparam prom_inst_33.INIT_RAM_2D = 256'hFFEFFEFFFFFFFFFFFFFFDF9FFAAFEBD7F9DFFD7AFFFBFFBFFD7BFFFE7FEBFFAD;
defparam prom_inst_33.INIT_RAM_2E = 256'hF77F5EBFFEBFFFFF5F5FFF9FFAFFF55FFF5FFE7FFD7FFFFFFFFFFFFFFFDFF7FF;
defparam prom_inst_33.INIT_RAM_2F = 256'hD7FF9FFF5FFFFFFFFFFF7FFFFFFFFFFFFFFF7FFFFFFFFFFFFFF7EBFE2BF9FAFE;
defparam prom_inst_33.INIT_RAM_30 = 256'h7F3FFFFFFFFFFFFFFFFAFFD0FFFEBFAF5FD7AFFFAFFFFFCFD7F5EFFEBFFE97FF;
defparam prom_inst_33.INIT_RAM_31 = 256'hF40FFC0BFFFFF3FDFD72FFAFFFA5FE05FFE7F817FFFFFFFFFFDFFFFEFFBFFFFF;
defparam prom_inst_33.INIT_RAM_32 = 256'hFAFEFDFFFFFFFFFFFFFFFFFFEFFFFFDF3FFFFFFFFFFFFFFFFEBFF6BFFFAFEA97;
defparam prom_inst_33.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFEFAFFEF7FFFBFAAFFDFFFF7EFFDFFCFEFFA1BFFBFFEF7FFF7F;
defparam prom_inst_33.INIT_RAM_34 = 256'hFFC0FFF5FF5FBFEFEFFEFFFADFE05FFEBF807FFFFFFFFFFEFFFFFFFFFFFFF81F;
defparam prom_inst_33.INIT_RAM_35 = 256'hFFAFFFFFFFFFFFBFFFFDFF7FFFFFFFFFFFFFFFFFFFFFFBEBFF4DFFFCFEA7FF60;
defparam prom_inst_33.INIT_RAM_36 = 256'hFFFFFFFFFFFEFAFFD37FFF3FA1FFE3FFFFFFFD7FD7EFFB1BFFFFFD97FFD7FFAF;
defparam prom_inst_33.INIT_RAM_37 = 256'hFFFF5FF5FBFEBAFFDFFF5AFFF9FFEBFFEBFFFFFFFFFFF7FFFFFFDFFFFFFFFFFF;
defparam prom_inst_33.INIT_RAM_38 = 256'hFFFFFFFFFFFDFFFFEFFFFFFFF80000FFFFFFFFFFFFBF3FEF5FFFDFF17FF8F7FF;
defparam prom_inst_33.INIT_RAM_39 = 256'hFFFFFFFFEFCFFAD7F3FFFDBBFEBD7FFFFFF7FF7EFFAF3FF7FFF6BFFE7FFAFFFA;
defparam prom_inst_33.INIT_RAM_3A = 256'hFFFFAFFFEFCFFD7FEFAFFFAFFFBFFEBFFFFFFFFFFFFFFFFBFEFFFFFDFFFF9FFF;
defparam prom_inst_33.INIT_RAM_3B = 256'hFFFFFFFFEFFFFFFFBFFFFF7FFFF9FFFFFFFFFFFBF3FFB5FD7AFF6EBFAF5FFF5F;
defparam prom_inst_33.INIT_RAM_3C = 256'hFFFFFEFD7F7F7FCCBFDBAFEBD7FBB7FFFFF1D7FAF7FF5FFAEBFFCBFFAFFFAFFF;
defparam prom_inst_33.INIT_RAM_3D = 256'hFD8DFEBD7FD7FFBAFE06FC1BF81BFFFFFFFFFFFBFFFFDFFFFFFFEFFFFFBFFFFF;
defparam prom_inst_33.INIT_RAM_3E = 256'hFFFFFFFFFFF7FDFFFFFBFFFFF7FFFFFFFFFFBF5FD79FEC6FF6EBFAFDFD0DFFFF;
defparam prom_inst_33.INIT_RAM_3F = 256'hFFEFD7FDEBFDF7FD7EFEBFFF7F7FFFFFB6FFAF5FF5FF7EBFBFBF7F7EFEFFFFFF;

pROM prom_inst_34 (
    .DO({prom_inst_34_dout_w[30:0],prom_inst_34_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_34.READ_MODE = 1'b1;
defparam prom_inst_34.BIT_WIDTH = 1;
defparam prom_inst_34.RESET_MODE = "SYNC";
defparam prom_inst_34.INIT_RAM_00 = 256'h3FE3CFFE7FC7CFE00FC03FC03FFFFFFFFFFFDFFFFFFFFFFFFEFFFFFE7FFFFFFF;
defparam prom_inst_34.INIT_RAM_01 = 256'hFFF7FFFFBFEFFFFFDFFFFFDFFFFFFFFFFBF1FCF9FF81FF1F3FCF9FC01FF9FFF0;
defparam prom_inst_34.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFBFFFFF7FFFFFBFFFFFFFFFE;
defparam prom_inst_34.INIT_RAM_04 = 256'hBFFFFFFFFFFFFDFFFFFF7FFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FDFFFFFBFFFFFDFFFFFFFFFEFFF;
defparam prom_inst_34.INIT_RAM_07 = 256'hFFDFF7FFFFEFFFFFFBFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFBFFFFFFFBFFFFFEFFFFFFFFFEFFFFFF;
defparam prom_inst_34.INIT_RAM_0A = 256'hFFBFFFFEFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFE;
defparam prom_inst_34.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFDFFFFFF7FFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_0D = 256'hFFFFF7FFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FD;
defparam prom_inst_34.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFBFFFFDFF7FFFFDFFFFFFBFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_10 = 256'hFF7FFFFFEFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_11 = 256'h3FE07F8FF07FFCF3FF80780F00FE7DF3CF3FCFC07FFFFFFFFFFFF7FFFF7FDFFF;
defparam prom_inst_34.INIT_RAM_12 = 256'hFFEFF7EFFFFFFFFFFFFDFFFFEFFBFFFFDFFFFFFBFFFFFFFFDFFCF3CF9C03CFFF;
defparam prom_inst_34.INIT_RAM_13 = 256'hFFFFFEFFFFFFFFF7FFBD7BFF7EF7FFBFF7EFFBFBEFFFBD7FFFEDFFDFDF9EBDFD;
defparam prom_inst_34.INIT_RAM_14 = 256'h0FFFFE85FFCF5FF8C78171C7EBEF5E35FB7C0BFFFFFFFFFFFFFFFFFBFEFFFFF7;
defparam prom_inst_34.INIT_RAM_15 = 256'hFFFAFFFFFFFFFFFFEFFFFF7FDFFFFDFFFFFFBFFFFFFFFFFFCF5D7FC0BD7FEDFF;
defparam prom_inst_34.INIT_RAM_16 = 256'hFFEFFFFFFFFEFFF7F75F781F5FFBFEDBFFDFACFFF3F7FF51FF5E23FAFFD78D7E;
defparam prom_inst_34.INIT_RAM_17 = 256'hC7E7BFFD7FFFF5FFFFEBFEBFF5F5DFABFFBFFFFFFFFFFFFBFFFFDFF7FFFF7FFF;
defparam prom_inst_34.INIT_RAM_18 = 256'hCFFFFFFFFFFFFF7FFFF7FDFFFFDFFFFFFBFFFFFFFFBFFD7DE7DFF5F7FEAFEF7F;
defparam prom_inst_34.INIT_RAM_19 = 256'hFFFFFFFFEFFF5EFAF7FD7DFFFBFBD7D2FFEBFF5FFFFF7FFFFEFFAFFD7EB7E4FF;
defparam prom_inst_34.INIT_RAM_1A = 256'hF2FFD7FFFFDFFFFFBFF3DF9FF7FD7FF3FFFFFFFFFFFFDFFFFEFFBFFFF7FFFFFE;
defparam prom_inst_34.INIT_RAM_1B = 256'hFFFFFFFFFFF7FFFFBFEFFFFDFFFFFFBFFFFFFFF7FFD7BEBDFFDEFFFDFEF5F5BF;
defparam prom_inst_34.INIT_RAM_1C = 256'hFFFFFDFFFDEFCF7C17BFFF5F5D7D5FF1BFFDEBFFEFF07FDFFCF5E7FDFF77C3FF;
defparam prom_inst_34.INIT_RAM_1D = 256'hFE7AFFFBFDFBF5FF3F7AFDFFDFEFDFFFFFFFFFFFFEFFFFEFFBFFFF7FFFFFEFFF;
defparam prom_inst_34.INIT_RAM_1E = 256'hFFFFFFFFBFFFFDFEFFFFBFFFFFFBFFFFFFFFFFFF7AF5DEFFEBFFE7F85F55FBDF;
defparam prom_inst_34.INIT_RAM_1F = 256'hFFBFFFBEBE57C1FAFFDAFBFFDF7DCFFF9FBFFEFF02FD7FD7DEBFDBF6BC17FFFF;
defparam prom_inst_34.INIT_RAM_20 = 256'hEFFFAFFEBF5FF5FFAFA2FDAF85FFFFFFFFFFFFEFFFFF7FBFFFEFFFFFFDFFFFFF;
defparam prom_inst_34.INIT_RAM_21 = 256'hFFFFFDFFFFEFCFFFFBFFFFFF7FFFFFFFEFFFEFEF97FF2EBFFEBEC7F5FF47FFEF;
defparam prom_inst_34.INIT_RAM_22 = 256'hFFFAF3E9FFEBCE7E3FAEFD0BD7FFFAFFFFEBFFFFF7FD7FEBEABD8FFF7FFFFFFF;
defparam prom_inst_34.INIT_RAM_23 = 256'hFEFFF7FDFFDEFAFFCF637FBFFFFFFFFFFFFE7FFFFBF7FFFDFFFFFF9FFFFFFFF7;
defparam prom_inst_34.INIT_RAM_24 = 256'h0FBFFFFF03FFFF7FFFFFEFFFFFFFFBFFFEBDFC7FFEF39F8DEBAF66F5E7FFBDFF;
defparam prom_inst_34.INIT_RAM_25 = 256'hFF7F5FFFFDE7FF7AEBDFFCFFFFFF7FFF3FFDFEFFE7AEBDF7DFDFEFFFFFFFFE00;
defparam prom_inst_34.INIT_RAM_26 = 256'hE0DFBF01F9AF5DF5EFFAFFFFFFFF8003FFFFFFE0FFFF3FFFFFF7FFFFFFFCFFFF;
defparam prom_inst_34.INIT_RAM_27 = 256'hFFFFF800001FFFFFFFFFFFFFFF7FFFF5BFFFFFBF59D7AEBEF5D75DFFF5BFFFDF;
defparam prom_inst_34.INIT_RAM_28 = 256'hFFFC0FD175EBAF3EFFE0DFFF8FFFF7F837EBC3BD1BF75D7AFEBFFFFFFFE00000;
defparam prom_inst_34.INIT_RAM_29 = 256'hFAF7EFBFFFD75FBFEFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFCFFFFFFFFBFFFFD8F;
defparam prom_inst_34.INIT_RAM_2A = 256'hFFFFFFFFFFFFFE7FFFFFFFDFFFFFB6FEFF7FFADD7CEBDFBEB97FFFBEFFFD7FFD;
defparam prom_inst_34.INIT_RAM_2B = 256'hC03F073F3CF3CFCF03FFF07FFF3F807F3C03F07CFBEFCFF3FFFFFFFFFFFFF7FF;
defparam prom_inst_34.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEFFFFFFFFFFF7FFFFFFFEFFFFFF07FCF;
defparam prom_inst_34.INIT_RAM_2D = 256'hFFFFFFFFFC1FFFFFFFE7FFFFFF3FFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF0000000000FFFFFFFFF3FFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_30 = 256'h07FFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFE000;
defparam prom_inst_34.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_33 = 256'hFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFF7FFFFC0000000000000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_3B = 256'hFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFBFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_34.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_35 (
    .DO({prom_inst_35_dout_w[30:0],prom_inst_35_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_35.READ_MODE = 1'b1;
defparam prom_inst_35.BIT_WIDTH = 1;
defparam prom_inst_35.RESET_MODE = "SYNC";
defparam prom_inst_35.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00F;
defparam prom_inst_35.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0007FF;
defparam prom_inst_35.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFF;
defparam prom_inst_35.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFF;
defparam prom_inst_35.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_12 = 256'hFFFFFFFFFFFFF80000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_15 = 256'hFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_18 = 256'hFFFFFFFC00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800003FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1B = 256'hFFFFE00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1E = 256'hFF000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_21 = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam prom_inst_35.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_24 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_35.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000F;
defparam prom_inst_35.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFF;
defparam prom_inst_35.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000003FFFFFF;
defparam prom_inst_35.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFF;
defparam prom_inst_35.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFC000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_35 = 256'hFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_38 = 256'hFFFFFFFFFE000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3B = 256'hFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3E = 256'hFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_35.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_36 (
    .DO({prom_inst_36_dout_w[30:0],prom_inst_36_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_36.READ_MODE = 1'b1;
defparam prom_inst_36.BIT_WIDTH = 1;
defparam prom_inst_36.RESET_MODE = "SYNC";
defparam prom_inst_36.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000003FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_01 = 256'hFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam prom_inst_36.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_07 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000;
defparam prom_inst_36.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000003F;
defparam prom_inst_36.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFF;
defparam prom_inst_36.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFF;
defparam prom_inst_36.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFF800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_18 = 256'hFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_1B = 256'hFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_1E = 256'hFFFFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_21 = 256'hFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_24 = 256'hF000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_27 = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam prom_inst_36.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_2A = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000;
defparam prom_inst_36.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FF;
defparam prom_inst_36.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFF;
defparam prom_inst_36.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFF000000FFFFFF800003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_33 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000;
defparam prom_inst_36.INIT_RAM_35 = 256'hFFFF800000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_36 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000;
defparam prom_inst_36.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFC000003FFFE0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_39 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFE00000000;
defparam prom_inst_36.INIT_RAM_3B = 256'hFFFFFFFFFFFE000007FFFFE0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_3D = 256'hFFFFEFFFFFFF7FFFFFFFFDFFFFFFFFFFFFFFFFFFFFC00000FFFFFC0000000001;
defparam prom_inst_36.INIT_RAM_3E = 256'hFFFFFFFFF000003FFFFF80000000003FFFFEFFFFFFFFFFF7FFFFFFFFFFFFFFFF;
defparam prom_inst_36.INIT_RAM_3F = 256'hFFBFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_37 (
    .DO({prom_inst_37_dout_w[30:0],prom_inst_37_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_37.READ_MODE = 1'b1;
defparam prom_inst_37.BIT_WIDTH = 1;
defparam prom_inst_37.RESET_MODE = "SYNC";
defparam prom_inst_37.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFC00000FFFFFE00000000003FF;
defparam prom_inst_37.INIT_RAM_01 = 256'hFFFFFF800001FFFFFE0000000000FFFFFFFFFFFF7FFF7FFF7FFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_02 = 256'hFFFFFFDFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_03 = 256'hFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007FFFFF80000000000FFFFF;
defparam prom_inst_37.INIT_RAM_04 = 256'hFFF800001FFFFFF00000000001FFFFFFFFFFF7FFF7FFFFFFFFFFFFFFFFFFFFF7;
defparam prom_inst_37.INIT_RAM_05 = 256'hFFFFFFFDFFFFFFFFFFFFFFFFFFFFFDFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFF0000000001FFF000003FFFFFE00000000003FFFFFFF;
defparam prom_inst_37.INIT_RAM_07 = 256'hC00000FFFFFF800000000007FFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_08 = 256'hEFFFDFFDEFFFFDFFFFEFFFFFFFFFFFDFFFFFFFFFFEFFFFFFFFFE0000000001FF;
defparam prom_inst_37.INIT_RAM_09 = 256'hFFFFFFFFBFFFFFFFFFFFFFF000007FF000003FFFFFF00000000001FFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_0A = 256'h0007FFFFFC00000000003FFFFFFFFFFBFFF7FFFFFF7FFFFFFBFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_0B = 256'hFDFFFFFFFFFFFFFFFFFFFFFEFFFFFFF7FFFFFFFFFF7FFFFFFFFFFC00000FFE00;
defparam prom_inst_37.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFF800003FF800001FFFFFF000000000007FFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_0D = 256'h7FFFFFE00000000001FFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFBFFFFFFDFF;
defparam prom_inst_37.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007FF00000;
defparam prom_inst_37.INIT_RAM_0F = 256'hFFFFFEFFFFFFFFFFFC00001FFC00000FFFFFF800000000003FFFFFFFFFFFFFDF;
defparam prom_inst_37.INIT_RAM_10 = 256'hFFFE000000000007FFFFFFFFFFFFF7FFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_11 = 256'hFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FF000003FF;
defparam prom_inst_37.INIT_RAM_12 = 256'hFFF7FFFFFFFFFFF00000FFE000007FFFFFC00000000001FFFFFFFFFFFFFDFFDF;
defparam prom_inst_37.INIT_RAM_13 = 256'hF000000000003FFFFFFBFFFFFF7FF7FFFFFFFFFFDFFFFFFFDFFFFFFEFFFFDFFE;
defparam prom_inst_37.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FF800001FFFFF;
defparam prom_inst_37.INIT_RAM_15 = 256'hFFFFFFFFFFFF80000FFE000007FFFFFC00000000000FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_16 = 256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFC00000FFFFFF00;
defparam prom_inst_37.INIT_RAM_18 = 256'hFFFFFFFFFC00007FF000003FFFFFC000000000007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_19 = 256'h0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFE00000FFFFFF00000;
defparam prom_inst_37.INIT_RAM_1B = 256'hFFFFFFE00003FF800001FFFFFC000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_1C = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000FFE000003FFFFE00000000;
defparam prom_inst_37.INIT_RAM_1E = 256'hFFFE00001FFC00000FFFFF8000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_1F = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00007FF000003FFFFE00000000000;
defparam prom_inst_37.INIT_RAM_21 = 256'hF00001FFC00000FFFFF8000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FF800001FFFFC0000000000003F;
defparam prom_inst_37.INIT_RAM_24 = 256'h000FFE000007FFFF0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam prom_inst_37.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FF800001FFFF80000000000001FFFF;
defparam prom_inst_37.INIT_RAM_27 = 256'h7FF000003FFFE00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_37.INIT_RAM_28 = 256'hFE0FFEFCFF7E7F807F007FC1FFE03FC03FDFFFC07FFEFF00FFFFFFFFFFF80000;
defparam prom_inst_37.INIT_RAM_29 = 256'hFBEFFFDFFFBFFF3FFFFFFFFFFE00001FFC00000FFFF80000000000001FEFF9F7;
defparam prom_inst_37.INIT_RAM_2A = 256'h000001FFFC00000000000003FBFF7DFFBDFFBE3FFFDFFF9FFCFFF7BFF9EFFE7F;
defparam prom_inst_37.INIT_RAM_2B = 256'h3FFF8FFBF7FFE7FF3FFBF7FCFBFF9FFE7BFFFFFFEFFFEFFFFFFFFFFFC00003FF;
defparam prom_inst_37.INIT_RAM_2C = 256'hFFFFFFFBFFFBFFFFFFFFFFF00000FFE000007FFE00000000000000FFFFEF7FCF;
defparam prom_inst_37.INIT_RAM_2D = 256'h001FFF000000000000003FFFFDDFF7EFFFE3FEFDFFFDFFCFFEFCFF3FFFF7FFDE;
defparam prom_inst_37.INIT_RAM_2E = 256'h78FFBF7FFF7FF3FFBFBFCFFFFDFFFBBFFFBFFFFFFEFFFFFFFFFFFC00003FF800;
defparam prom_inst_37.INIT_RAM_2F = 256'hEFFFFFFFBFFFFFFFFFFF800007FE000003FF800000000000000FF7FFF7FFFDFF;
defparam prom_inst_37.INIT_RAM_30 = 256'hFFC000000000000001FDFFEFFFFF7FDCBFEFDFFFDFFCFFFFEFFBF7FF7FFF6FFF;
defparam prom_inst_37.INIT_RAM_31 = 256'hFBF3FFF7FF3FFFFBFEFDFFDFFFDBFFFBFFFFFFEFFFFFFFFFFFE00001FFC00000;
defparam prom_inst_37.INIT_RAM_32 = 256'hFDFF03FFFFFFFFFFF800003FF000003FC0000000000000007F7FF97FFFDFF76F;
defparam prom_inst_37.INIT_RAM_33 = 256'h000000000000001FDFFF0FFFF7FDD9FE00FF81FFEFFFFF7FDE7FF7FFF0FF80FF;
defparam prom_inst_37.INIT_RAM_34 = 256'h3FFF3FFBFFBFDFF01FFDFFFD3FFFBFFF7FFFFFFFFFFFFFFF00000FFC000007E0;
defparam prom_inst_37.INIT_RAM_35 = 256'hFFDFFFFFFFFFFFC00003FF800000000000000000000007F7FFB3FFFFFF7E7F9F;
defparam prom_inst_37.INIT_RAM_36 = 256'h000000000001FDFFECFFFFFFDF9FFFCFFFCFFEFFEFF7FCE7FF3FFE6FFFEFFFDF;
defparam prom_inst_37.INIT_RAM_37 = 256'hF3FFBFFBFDFF7DFFEFFFBDFFFFFFF7FFF7FFFFFFFFFFF800007FE00000000000;
defparam prom_inst_37.INIT_RAM_38 = 256'hFFFFFFFFFFFE00001FF8000007FFFF0000000000007FFFF3BFFFEFFEE7FFFBFF;
defparam prom_inst_37.INIT_RAM_39 = 256'h000000001FFFFDEFFFF3FE7DFF7EFFFCFFEFFEFF7FDFFFFBFFCF7FFFFFFDFFFD;
defparam prom_inst_37.INIT_RAM_3A = 256'hF9FFDF9FF7FFFEFFF3DFFFDFFF7FFF7FFFFFFFFFFF800007FF000003FFFFE000;
defparam prom_inst_37.INIT_RAM_3B = 256'hFFFFFFFFF00000FFC00000FFFFFE000000000007FFFE7BFEFDFF9F7FDFBFFFBF;
defparam prom_inst_37.INIT_RAM_3C = 256'h000001FEFF9EFFBF7FE7DFF7EFFFCFFE7FFFEFFDFBFFBFFDF7FFF7FFDFFFDFFF;
defparam prom_inst_37.INIT_RAM_3D = 256'hFE73FF7EFFEFFE7DFFF9FFE7FFE7FFFFFFFFFFFC00003FF000001FFFFFC00000;
defparam prom_inst_37.INIT_RAM_3E = 256'hFFFFFF00000FFE000007FFFFF800000000007FBFEFFFF39FF9F7FDFBFEF3FF9F;
defparam prom_inst_37.INIT_RAM_3F = 256'h001FEFF3F7FE0FFEFDFF7E7F80FFE7FFC9FFDFBFFBFF9F7FC07F80FF01FFFFFF;

pROM prom_inst_38 (
    .DO({prom_inst_38_dout_w[30:0],prom_inst_38_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_38.READ_MODE = 1'b1;
defparam prom_inst_38.BIT_WIDTH = 1;
defparam prom_inst_38.RESET_MODE = "SYNC";
defparam prom_inst_38.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FF800001FFFFFF80000000;
defparam prom_inst_38.INIT_RAM_01 = 256'hFFF800007FF000003FFFFFE00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFC00000FFFFFFC0000000001;
defparam prom_inst_38.INIT_RAM_04 = 256'hC00003FF000003FFFFFF80000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFE000007FFFFFE0000000001FFF;
defparam prom_inst_38.INIT_RAM_07 = 256'h003FF800001FFFFFFC0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam prom_inst_38.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FE000007FFFFFF0000000001FFFFFF;
defparam prom_inst_38.INIT_RAM_0A = 256'hFFC00001FFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001;
defparam prom_inst_38.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF800003FF000003FFFFFF8000000001FFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0D = 256'h00000FFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFE;
defparam prom_inst_38.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFC00003FF800003FFFFFFC000000001FFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_10 = 256'h00FFFFFFF000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000FFE000;
defparam prom_inst_38.INIT_RAM_12 = 256'hCFF3F81FFFFFFFFFFFFE00001FFC00003FFFFFFC000000003FFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_13 = 256'hFFFFFF000000000FFF7EF7E781FBFFCFF81FE7FC1FFF7EFFE01E03E03FFF7EF3;
defparam prom_inst_38.INIT_RAM_14 = 256'hF3F8FF7BFFFFBFFF3FFEFE3FF7DFBFFBFCFFF7FFFFFFFFFFFF800007FF00000F;
defparam prom_inst_38.INIT_RAM_15 = 256'h1FFDFFFFFFFFFFFFF00000FFE00003FFFFFFC000000003FFFFBEF9FF7EFFF3FC;
defparam prom_inst_38.INIT_RAM_16 = 256'hFFF000000001FFFBEFBEFFEFBFFC7F3CFE3FDF7FFFEFFFEFFFBFDFFDF3EFFEFF;
defparam prom_inst_38.INIT_RAM_17 = 256'hBFFFDFFEF9FFFBFFE7F7FF7CFBFBBFD7FF7FFFFFFFFFFFFC00003FF80000FFFF;
defparam prom_inst_38.INIT_RAM_18 = 256'hFFFFFFFFFFFFFF80000FFE00003FFFFFFC000000007FFEFBFFBFFBEFFF5FDFBF;
defparam prom_inst_38.INIT_RAM_19 = 256'h000000001FFFBF7DEFFEFBFF97F7EFEDFFF7FFBE7FFEFFF9FDFFDF3EFF6FFFFF;
defparam prom_inst_38.INIT_RAM_1A = 256'hFDFFEF9FFFBFFE7F7FFFEFFFC9FBBFFFFFFFFFFFFFFFE00001FFC0000FFFFFFF;
defparam prom_inst_38.INIT_RAM_1B = 256'hFFFFFFFFFFF800007FF00003FFFFFFC00000000FFFEFDF7BFFBF7FE6FDFBFB7F;
defparam prom_inst_38.INIT_RAM_1C = 256'h000003FFFBF7FEFFEFDFF9BFBEFEEFFE7FFBF7FFF7FF9FEFFFFBFFF27EEFFCFF;
defparam prom_inst_38.INIT_RAM_1D = 256'hFFFDFFFDFE07FBFFFEFDFE1FB9F03FFFFFFFFFFFFF00001FFC0000FFFFFFF000;
defparam prom_inst_38.INIT_RAM_1E = 256'hFFFFFFFFC00003FF00007FFFFFFC00000000FFFEFDFBBF01F7FE7FE7BFBBFC3F;
defparam prom_inst_38.INIT_RAM_1F = 256'h007FFFDF7FEFFE7DFFBDFC07EEFE3FFFFF7FFF7FFDFEFFEFBF7F27EF7FEFFFFF;
defparam prom_inst_38.INIT_RAM_20 = 256'hDFFFDFFF7FBFFBE7DFDDFBDFFBFFFFFFFFFFFFF00000FFC0001FFFFFFE000000;
defparam prom_inst_38.INIT_RAM_21 = 256'hFFFFFE00001FF00007FFFFFF800000001FFFF7DFFBFFDF7FE77F39FB9FBFFFF7;
defparam prom_inst_38.INIT_RAM_22 = 256'hFFFDFFF6FFF7FFF9CFDF7EF7EFFFFDF3FFF7FFCFEFFEF9F7F77E73FEFFFFFFFF;
defparam prom_inst_38.INIT_RAM_23 = 256'hFDFFFBFBFFBF7DF9FF9CFFDFFFFFFFFFFFFF800007F80003FFFFFFE00000000F;
defparam prom_inst_38.INIT_RAM_24 = 256'hF0400000FC0000FFFFFFF000000007FFFF7EFFBFFDFFFE73F7DF99FBFFFF7EFF;
defparam prom_inst_38.INIT_RAM_25 = 256'hCFBFAFFF3EFF80FDF7E03FF9FFCFBFFFFFFEFF7FFFDF7E7BE03FF7FFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_26 = 256'hFF3FDFFFF7DFBEFBF7FDFFFFFFFFFFFC0000001F0000FFFFFFF800000003FFFF;
defparam prom_inst_38.INIT_RAM_27 = 256'h000007FFFFFFFFFFFC00000000FFFFFBCFE3FFCFBFEFDF7DFBEFBE7FFBCFFFEF;
defparam prom_inst_38.INIT_RAM_28 = 256'hF8FFF3EEFBF7DFFDF9FF3FFE73FFFBFFCFF7FC7EE7CFBEFDFF7FFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_29 = 256'hFDF81FC1F3EFBF7FDFFFFFFFFFFFFFC00001FFFFFFFFFFFF000000007FFFFE73;
defparam prom_inst_38.INIT_RAM_2A = 256'h007FFFFFFFFFFF800000003FFFFFC9FF3F80FD3EFFF7EF7F7E8FFFC1FFFEFE03;
defparam prom_inst_38.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800;
defparam prom_inst_38.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFF800000001FFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2D = 256'hFFFFFFFFFFE00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800003;
defparam prom_inst_38.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFF000000000FFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_30 = 256'hF80000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00001FFF;
defparam prom_inst_38.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFF00000000000000000000003FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_33 = 256'h00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000;
defparam prom_inst_38.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFF800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FFFFFFFFF;
defparam prom_inst_38.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3B = 256'hFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3E = 256'hFFFFFFFFFFE00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_38.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_39 (
    .DO({prom_inst_39_dout_w[30:0],prom_inst_39_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_39.READ_MODE = 1'b1;
defparam prom_inst_39.BIT_WIDTH = 1;
defparam prom_inst_39.RESET_MODE = "SYNC";
defparam prom_inst_39.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800005FFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_01 = 256'hFFFFFFFE000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800001FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_04 = 256'hFFFFEC00023FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000007FFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_07 = 256'hFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80001FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0A = 256'h00002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA;
defparam prom_inst_39.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800003FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0D = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB000;
defparam prom_inst_39.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF400005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007;
defparam prom_inst_39.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE00005FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000FFFF;
defparam prom_inst_39.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFF;
defparam prom_inst_39.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA00007FFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFE80001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00001FFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1E = 256'hFFFFFFFFFFFFE80000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD000037FFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_21 = 256'hFFFFFFFFFF000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD000017FFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_24 = 256'hFFFFFFFE00004FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000BFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_27 = 256'hFFFFA00002FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF900009FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2A = 256'hFC000017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2D = 256'h0001BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8;
defparam prom_inst_39.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_30 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000;
defparam prom_inst_39.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFD000017FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD00001F;
defparam prom_inst_39.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFD00000BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFF;
defparam prom_inst_39.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFE800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000017FFFFFF;
defparam prom_inst_39.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFC00027FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD00000FFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFF800012FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_39.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_40 (
    .DO({prom_inst_40_dout_w[30:0],prom_inst_40_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_40.READ_MODE = 1'b1;
defparam prom_inst_40.BIT_WIDTH = 1;
defparam prom_inst_40.RESET_MODE = "SYNC";
defparam prom_inst_40.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFDFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFCFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_04 = 256'hFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_07 = 256'hFF7FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0A = 256'hFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFF;
defparam prom_inst_40.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFE7;
defparam prom_inst_40.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFF;
defparam prom_inst_40.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFF9FFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFBFFFFFF;
defparam prom_inst_40.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFCFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1E = 256'hFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_21 = 256'hFFFFFFFFFF3FFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_24 = 256'hFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFBFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_27 = 256'hFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2A = 256'hFCFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_40.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_30 = 256'hFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFDF;
defparam prom_inst_40.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFEFFFF;
defparam prom_inst_40.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFF;
defparam prom_inst_40.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF7FFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_40.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_41 (
    .DO({prom_inst_41_dout_w[30:0],prom_inst_41_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_41.READ_MODE = 1'b1;
defparam prom_inst_41.BIT_WIDTH = 1;
defparam prom_inst_41.RESET_MODE = "SYNC";
defparam prom_inst_41.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_01 = 256'hFFFFFFFEFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_07 = 256'hFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0A = 256'hFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB;
defparam prom_inst_41.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0D = 256'hFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFF;
defparam prom_inst_41.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF;
defparam prom_inst_41.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FFF;
defparam prom_inst_41.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFDFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFBFFFFFF;
defparam prom_inst_41.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFDFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFDFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFEFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFDFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1E = 256'hFFFFFFFFFFFFF7FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_21 = 256'hFFFFFFFFFFBFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_24 = 256'hFFFFFFFBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_27 = 256'hFFFFDFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFBFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2A = 256'hFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_30 = 256'hFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF;
defparam prom_inst_41.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFF;
defparam prom_inst_41.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFF7FFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFEFFFFFFF;
defparam prom_inst_41.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF7FFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_41.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_42 (
    .DO({prom_inst_42_dout_w[30:0],prom_inst_42_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_4),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_42.READ_MODE = 1'b1;
defparam prom_inst_42.BIT_WIDTH = 1;
defparam prom_inst_42.RESET_MODE = "SYNC";
defparam prom_inst_42.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_01 = 256'hFFFFFFFF00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_04 = 256'hFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_07 = 256'hFF800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0A = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_42.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0D = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000;
defparam prom_inst_42.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001F;
defparam prom_inst_42.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFF;
defparam prom_inst_42.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFE00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFF;
defparam prom_inst_42.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00003FFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1E = 256'hFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_21 = 256'hFFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_24 = 256'hFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_27 = 256'hFFFFE00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2A = 256'hFF00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2D = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam prom_inst_42.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_30 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam prom_inst_42.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003F;
defparam prom_inst_42.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00001FFFF;
defparam prom_inst_42.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFF800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00001FFFFFFF;
defparam prom_inst_42.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFF800003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000FFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_42.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_43 (
    .DO({prom_inst_43_dout_w[29:0],prom_inst_43_dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_43.READ_MODE = 1'b1;
defparam prom_inst_43.BIT_WIDTH = 2;
defparam prom_inst_43.RESET_MODE = "SYNC";
defparam prom_inst_43.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE2AAAAAAABACFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFF7AAAAAAAAA97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFDAAAAAAAAAB3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFDEBAAAAAAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_0F = 256'hFFFFFFFFFFFFFF7AAAAAAAAA1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_12 = 256'hFFFFFFFFFFF3ABAAAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_15 = 256'hFFFFFFFF9EAAAAAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_18 = 256'hFFFFFFFAAAAAAAA83FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1B = 256'hFFE7AAAAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1E = 256'hCEAAAAAAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_21 = 256'hAAAAAAA0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9EA;
defparam prom_inst_43.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_24 = 256'hAAAAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3AAAA;
defparam prom_inst_43.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_27 = 256'hA9BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBAAAAAAA;
defparam prom_inst_43.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5EAAAAAAA83;
defparam prom_inst_43.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAABBFFF;
defparam prom_inst_43.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBAAAAAAAB6FFFFFF;
defparam prom_inst_43.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0EAAAAAAA0FFFFFFFFF;
defparam prom_inst_43.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAAAAAAADFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE8AAAAAAA87FFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9EAAAAAABFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_43.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_44 (
    .DO({prom_inst_44_dout_w[29:0],prom_inst_44_dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_6),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_44.READ_MODE = 1'b1;
defparam prom_inst_44.BIT_WIDTH = 2;
defparam prom_inst_44.RESET_MODE = "SYNC";
defparam prom_inst_44.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF95555555557FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF95555555556FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFD5555555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFE5555555555FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFF5555555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_0F = 256'hFFFFFFFFFFFFFF9555555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_12 = 256'hFFFFFFFFFFFD5555555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_15 = 256'hFFFFFFFFE5555555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_18 = 256'hFFFFFE5555555556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1B = 256'hFFF9555555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1E = 256'hA555555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_21 = 256'h5555555BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE55;
defparam prom_inst_44.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_24 = 256'h55556FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF95555;
defparam prom_inst_44.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_27 = 256'h56FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF95555555;
defparam prom_inst_44.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE555555556F;
defparam prom_inst_44.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE555555555BFFF;
defparam prom_inst_44.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF955555555BFFFFFF;
defparam prom_inst_44.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE55555555BFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE555555556FFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA55555556FFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE55555555BFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_44.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_45 (
    .DO({prom_inst_45_dout_w[27:0],prom_inst_45_dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_8),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_45.READ_MODE = 1'b1;
defparam prom_inst_45.BIT_WIDTH = 4;
defparam prom_inst_45.RESET_MODE = "SYNC";
defparam prom_inst_45.INIT_RAM_00 = 256'hFFFFFDA7666666666666679FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_06 = 256'hC8766666666666668DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0C = 256'h66666666667BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD9666;
defparam prom_inst_45.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_12 = 256'h666679FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC986666666;
defparam prom_inst_45.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_18 = 256'hDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA7666666666667;
defparam prom_inst_45.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDB987666666667AFFFFF;
defparam prom_inst_45.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDA87777777778FFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDCBBA998899AFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDCBA99ABCEFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_45.INIT_RAM_36 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_5 (
  .Q(dff_q_5),
  .D(dff_q_4),
  .CLK(clk),
  .CE(oce)
);
DFFE dff_inst_6 (
  .Q(dff_q_6),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_7 (
  .Q(dff_q_7),
  .D(dff_q_6),
  .CLK(clk),
  .CE(oce)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(prom_inst_20_dout[0]),
  .I1(prom_inst_22_dout[0]),
  .S0(dff_q_7)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(prom_inst_16_dout[0]),
  .I1(mux_o_12),
  .S0(dff_q_5)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_13),
  .I1(mux_o_14),
  .S0(dff_q_3)
);
MUX2 mux_inst_18 (
  .O(dout[0]),
  .I0(mux_o_16),
  .I1(mux_o_15),
  .S0(dff_q_1)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(prom_inst_20_dout[1]),
  .I1(prom_inst_22_dout[1]),
  .S0(dff_q_7)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(prom_inst_4_dout[1]),
  .I1(prom_inst_5_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(prom_inst_6_dout[1]),
  .I1(prom_inst_7_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(prom_inst_17_dout[1]),
  .I1(mux_o_31),
  .S0(dff_q_5)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_3)
);
MUX2 mux_inst_37 (
  .O(dout[1]),
  .I0(mux_o_35),
  .I1(mux_o_34),
  .S0(dff_q_1)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(prom_inst_21_dout[2]),
  .I1(prom_inst_22_dout[2]),
  .S0(dff_q_7)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(prom_inst_8_dout[2]),
  .I1(prom_inst_9_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(prom_inst_10_dout[2]),
  .I1(prom_inst_11_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(prom_inst_18_dout[2]),
  .I1(mux_o_50),
  .S0(dff_q_5)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_3)
);
MUX2 mux_inst_56 (
  .O(dout[2]),
  .I0(mux_o_54),
  .I1(mux_o_53),
  .S0(dff_q_1)
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(prom_inst_21_dout[3]),
  .I1(prom_inst_22_dout[3]),
  .S0(dff_q_7)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(prom_inst_12_dout[3]),
  .I1(prom_inst_13_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(prom_inst_14_dout[3]),
  .I1(prom_inst_15_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(prom_inst_19_dout[3]),
  .I1(mux_o_69),
  .S0(dff_q_5)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_3)
);
MUX2 mux_inst_75 (
  .O(dout[3]),
  .I0(mux_o_73),
  .I1(mux_o_72),
  .S0(dff_q_1)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(prom_inst_43_dout[4]),
  .I1(prom_inst_45_dout[4]),
  .S0(dff_q_7)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(prom_inst_23_dout[4]),
  .I1(prom_inst_24_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(prom_inst_25_dout[4]),
  .I1(prom_inst_26_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(prom_inst_39_dout[4]),
  .I1(mux_o_88),
  .S0(dff_q_5)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_89),
  .I1(mux_o_90),
  .S0(dff_q_3)
);
MUX2 mux_inst_94 (
  .O(dout[4]),
  .I0(mux_o_92),
  .I1(mux_o_91),
  .S0(dff_q_1)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(prom_inst_43_dout[5]),
  .I1(prom_inst_45_dout[5]),
  .S0(dff_q_7)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(prom_inst_27_dout[5]),
  .I1(prom_inst_28_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(prom_inst_29_dout[5]),
  .I1(prom_inst_30_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(prom_inst_40_dout[5]),
  .I1(mux_o_107),
  .S0(dff_q_5)
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(mux_o_108),
  .I1(mux_o_109),
  .S0(dff_q_3)
);
MUX2 mux_inst_113 (
  .O(dout[5]),
  .I0(mux_o_111),
  .I1(mux_o_110),
  .S0(dff_q_1)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(prom_inst_44_dout[6]),
  .I1(prom_inst_45_dout[6]),
  .S0(dff_q_7)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(prom_inst_31_dout[6]),
  .I1(prom_inst_32_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(prom_inst_33_dout[6]),
  .I1(prom_inst_34_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(prom_inst_41_dout[6]),
  .I1(mux_o_126),
  .S0(dff_q_5)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_127),
  .I1(mux_o_128),
  .S0(dff_q_3)
);
MUX2 mux_inst_132 (
  .O(dout[6]),
  .I0(mux_o_130),
  .I1(mux_o_129),
  .S0(dff_q_1)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(prom_inst_44_dout[7]),
  .I1(prom_inst_45_dout[7]),
  .S0(dff_q_7)
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(prom_inst_35_dout[7]),
  .I1(prom_inst_36_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(prom_inst_37_dout[7]),
  .I1(prom_inst_38_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(prom_inst_42_dout[7]),
  .I1(mux_o_145),
  .S0(dff_q_5)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(dff_q_3)
);
MUX2 mux_inst_151 (
  .O(dout[7]),
  .I0(mux_o_149),
  .I1(mux_o_148),
  .S0(dff_q_1)
);
endmodule //Gowin_pROM1
