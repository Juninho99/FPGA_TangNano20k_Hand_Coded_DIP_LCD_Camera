//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Tue Sep 05 14:35:08 2023

module Gowin_SDPB4 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);//gaussian_blur_5x5 - new

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [14:0] ada;
input [7:0] din;
input [14:0] adb;

wire lut_f_0;
wire lut_f_1;
wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [1:1] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [2:2] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [3:3] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [4:4] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [5:5] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [6:6] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [7:7] sdpb_inst_7_dout;
wire [23:0] sdpb_inst_8_dout_w;
wire [7:0] sdpb_inst_8_dout;
wire dff_q_0;
wire dff_q_1;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_0.INIT = 16'h0100;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_1.INIT = 16'h0100;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b1;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h777C3F10560BD618F9B39A9394FB7891D7B7BA203B00F8372CFD8FB585FB6A58;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hE79E03253EBE8088CA09797A16130109E165D428DF1DBAAE1BB97717B8638A1F;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h0B28EEC549F828E6AB0CCF2FB13143CB700182924F4F6442470606CD3A69B22E;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h3DB6E14F047FB08C115F5108FF2A48CDEA11C21D9E29F05C1E5550CB9C5C03FA;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hD00B26858F39BE7DB2A3340A5D887C05A24B5DD7E5A0CCECC104FADA5CD71E33;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hE4EC5D580D57DC830B168040044DA7400AC5DB4051840E5F8BA12C1E2D52E6D3;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h536206224BDC89AA7D19DEAFAEC379F77FB3E30B7115E820D21E34E6C1960F6C;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h5A4D9C6F16D52330FC5B86605D9407ADEC46CB8DEB81BBFCD9F93F7B427E7D7C;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h8A0CC1038FEA51C8556D47E9491DD17F5FAC7FFD9E30F0DFC07BF99BFB15EC23;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hAE7E864DE63C5348A7F24C09299446DEFFD4BBAE43F873E0376FD073C832662E;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h08E3EB2BBDCA68E12552A87F744EAF428D30C9CA369DD9148016FFFF8D897C2C;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h1B3CD40851B6D2D2AFBFBB827FDBDFEFFE9C58D33C5D7FD499309636E82F6925;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h63179E3B3F3DB5893FEC0013F73139D36101D84CEECC0ADE8D558C215104EDF0;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h054BFCC22B1ED36C80B57C92E8481DFD6B75500CAD75FEB8BBF597F2965554ED;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h7845C57578B9B4B885DEC4E091B5D33DE2D54F47E55E53BB0DBED559FE116586;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h9C2A2065203D91F2A7B28927652FE840DFFFCBF9DD883E19DB839B14E50FDAA9;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hA6E0BCEFC0EF8C5AA6EC06BCCABADAFC1154D803BBC1F20AACEFC2B8F1B8F31C;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h681103986673820D0D15F7E91A9F1B68ED90C40FD6C6B9CEDF4C9C9E5973E97C;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hBFCA7F51BCE32A4CD4DA52328B3EF8A401C0C94378BBB33EF2D8B0F046375EB4;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h66E2E247DF919E7F2DA2D6D77BD69EB096D6D106C0811A3457067904550080B4;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h094F9D9E06BB52F053067CEE45A0389F0DB5C8FD3CEF0E8FE604CB5F64764E69;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hF3BC247BF476198EDDE1FF0333B6AD83CCCC076C4B5985715F912A90CED49C3D;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h12D3F66CF6801204ABABC24F715810F4AD08EFCCB394AF8F945312E174BE9C8F;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hDC6515E23A2BBC2BF55C680DFFE7D74C55439C684402F8E9A95C1658A84C855D;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hD07F7C4C9E36272F1F2422FB702AC017146F7C6149723259D2B39E3167A8076E;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h1E0773AF38CDF3DFD8B89382FB947AEFE52BA70C09492ED4C05B49EE5EF50024;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hD4BDD072DDE02166340E96D4A2CBC2BFA6DFB45102D0B7CC542828DCB678181F;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h23CC75C12C6918F9A38F323B4A8F1B6F44EB4B44EEF8FF457C3F8292CDC47B0F;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h13E426A89DF69B410B91003A0FB031DFC0476FFC1D51993AFB1A2F52D2EF891A;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h084ADE4D816AF827803699BEEAD39C175386EF6A8AAEC0F9904FA4BCE90F1FCB;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h126935A9B9FC541077630C6B282A1B0737BA05AFB72C274FCB8159642D6DFD80;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h58F883B9F7BE877FE08D5865CD624A2503FD9ED7A08F9378601078712D548810;
defparam sdpb_inst_0.INIT_RAM_20 = 256'hC52A62213634BDBB2771CF9E9CC5F094690AFFD34B427F9DAF58001A1B2E2800;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h3E7ED9C4961AA6F4C7C9725E9E656B51089C532490584778145C3C6B46E40DC6;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0F8080B4023C55F06CE28DC7C5F1C0EF3756FD66476DFD606A6C5C3282A05BE6;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h5FF282E425FF2B5D7B9608785B42C03309BE4C6D9BB94C01377CDF4B5AF105C9;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h04D336A4CFBABEC013B0CDDB38BFC29BF6D801FF69ACD9D48044997D4AD3E450;
defparam sdpb_inst_0.INIT_RAM_25 = 256'hB60D0378DA117FFABD9C7DC3D87CB5FEC6C5A0CD24B8C143288B20B81EF0BABB;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h9BA6E43D09EC3700C4B35982FD081FFC229EF34FBC2E88B7BAB6C9136B023E3D;
defparam sdpb_inst_0.INIT_RAM_27 = 256'hF433ED2DE6F70BC9664587BFBFC20BC6282A570801F80BE29EBF65914C786439;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h8B9F10BC055338E79B681DE009FBBFBD6130C26ECF3AEF6421F4507B662F3F36;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h0FE7AF1BFF7ACB4ACD893EE73C77E3B7075F396437FA90E6BA9CDEB2BF6DB039;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0E2AFEA87FC0B802A0E148FC553347D10176E4937CFCFEF8D8400DECB3BF4DB7;
defparam sdpb_inst_0.INIT_RAM_2B = 256'hE93E6A7910F42AD9D09D7F941B4B72CF51408C14CAD4B78969B4D8CB4B0C5384;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h88CB93C7776BF96A2B7EBBFBED5F35AA6E9CC7939B10B002E13EF3CFAA11378D;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h3969B1FB1666A81D408DC40A928151D370953A5AF441C06E1C15BEF0200E24B8;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h6D50D3FB3D9258D9726F8F1A391F7E91AF46C5A7A65C2E5D8087FFDF832F42FE;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h51D51D61DC09436665555AE2742D62E575C2846DE7027AD8449C037482064472;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h4E27C5A02DFE41A0AC9B02C2EACDA7C72AE5E209694AC10E38EAF884862913EC;
defparam sdpb_inst_0.INIT_RAM_31 = 256'hA6F9A90B3143FF7DEC3B564755B7A566C36CB3149C9AC8FABF548D2FF0503AF0;
defparam sdpb_inst_0.INIT_RAM_32 = 256'hCB46F5F8E5D50F56D58A3E7F38ACD9967F46DC136130A558360C222FBA5FA797;
defparam sdpb_inst_0.INIT_RAM_33 = 256'hE1A8165FE2BBBC82DEBB33CBF9E69A88E21E6AEEC12B0723E7FBC8829C3AD9D4;
defparam sdpb_inst_0.INIT_RAM_34 = 256'hB000038543220B5224E4BBF5574C25FCFD6AB2F2ADCC49E929EDC55F120824E8;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h11FC334AEDA90EA164E1625F76FF0973DEB10D5F003DEE8CD3FEE612BDE76364;
defparam sdpb_inst_0.INIT_RAM_36 = 256'hEF2B18D9FB4FE28B63A693DC35C1717F44F259995D1C9D763F1E3644C6FC1AE0;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h1D1ABDDDCC127FF3B3EE2A6EBBF5F5047B83185FF8D3D6D90E10962146612E85;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h9CAEDD0914109EC40E877189645F90DB61DE491CFCC38E9B019F657156125466;
defparam sdpb_inst_0.INIT_RAM_39 = 256'hFAF898556A208034ADEF319B167D73757E98445E4B6C15C4ED86472FFE96D6AE;
defparam sdpb_inst_0.INIT_RAM_3A = 256'hB3556906AF716BD9F6E8D401BC9DDE5C87DE16AE45C1E51FBD7C6EB40DB7419F;
defparam sdpb_inst_0.INIT_RAM_3B = 256'hAEDE4CC32891C70BF6F4B79D4CFBB9B879A848A68DF327F7F03AB203D0A42C06;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h421B90E74F009495302677B90D9A15947E81BCED1168A62ACDABF3A2D291D1C1;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h9658AB7F114C5CC93840D4B980064CE6A9AE97B13C8BB5E444D96255010E89B6;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h2EA92EA1DC3B5EE2947627BBD0A138D462AF2C9AC7C8EB80962FFD2ED20AA447;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h804001319C868203A0CFBB2BDF5FCA46A49F7B952A12B9E605655AE2485F3851;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b1;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h5FFD2C5077CF8000F9EFDC99F506786FD0004DC0DCFFFFB33CFDBFE004FAFD56;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h0001FB00FE400FF7200D7BFA10010119F688062BF4DCA181EB23FD00F39C0A7F;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h0800010448FFD7080B0205924F70BDC002D27D124E470008230607BEC02B9FBF;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h827FE0BF007CFDC4117F5000000028CDFDFE20150E40079C01D401EEBFA003FA;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h000B20018F79FF8200201365DC07FC0EEE7EFFD7EDA008000204F3FFE2211500;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h1BFC42F87133C5B0FEEF8000000007FBFFFA24880A7FFE507FA17D63EB7FFED0;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h25600602EFDFFDC5906625FFA03B6F2DC2527CFFF0076001801E37FFFECA8803;
defparam sdpb_inst_1.INIT_RAM_07 = 256'hFA483CF71AA7D90003D059D710000FFDFFFF7462157FB8133CDEC2ECA3419D00;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h3C63E003AFFB5FFFBE92FFE806FB981880FDFE05235C4420007BFDFFFFCA42DF;
defparam sdpb_inst_1.INIT_RAM_09 = 256'hADA17A3D05F2FEC79603A39B160046FFFFFFDD31FDFC001FDEA2BE0ECFF164AF;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h3564326EBFFE6DFECA6FA0008B9690E086F7BBC83E474BE4841EF7FEDAF603EC;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h00820E3DBE03C141FFB0F1CA00005FEFFE1EE63FB4480029769E4E2A681F6997;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h3F80603B7F7DBFD677CE000806F3BCECD524878F11B1D02008558C3BF7CB79F0;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h880D7F64AF8252E876153486070A1DFD6B7EACFEAD7000AB53961AC6CE32ECF8;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h04C00577F8B9BE4FFDDFF5C056DD88757D4B9BD3E65170040FBED55FE3F5A7C6;
defparam sdpb_inst_1.INIT_RAM_0F = 256'hD3DFFAE5C9768315BCAE32D1622FFC40FF9077FBF690336B2ED9B63C3303DEAD;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hF9AABBFFE06EE2BEFF7A30F1A7E46B56C87B68B5E324260BAEEF42AE0FFEFE0D;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h65C1EDF890B7A922401264EEFFDF5B68FDC7EBE54F173D047B3E045ABB024DAA;
defparam sdpb_inst_1.INIT_RAM_12 = 256'hC071FF71E9FD97B72438528EC8C383017A8A26A61AD40C3E7EFB3A95B5C84372;
defparam sdpb_inst_1.INIT_RAM_13 = 256'hEDB7DE47657F07010F5BE017A5F69EB1F4292EA810171D0FC753579772EF3505;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h09F87D9E07D91C8F41FBC7438D529DE73EA04F278253147FE5456D109A882347;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h85CC39555C1EB0F35F65011D0FB70D9DA030077875123943ADA4E265C888B490;
defparam sdpb_inst_1.INIT_RAM_16 = 256'hE84FFE6EFD83820F4DFA2CC1FAA54BCA25A5160F0827747F9C579A1624BD1090;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h878F2926059079C790E4AC447FEFC79E240366B398F463E26B3E671902793ED1;
defparam sdpb_inst_1.INIT_RAM_18 = 256'hA5FF7C0E980807C8B9A3FE870FD9C3FD25E4FEB14A2A4FF9D23C900278CDE35E;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h05F88F81F8F025DF6F82B0DFFF1475804175FCC01DDF0115202FF2683EE3F8C2;
defparam sdpb_inst_1.INIT_RAM_1A = 256'hCEFDD07DC200264B3E1E71DFFEC03FBF202FB9624E2477CCDDDC128D456920F9;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h03C8023FAC682FFE354A25FBE88FF8004452400CB23CFDC483FF8083EDAA8E91;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hB764E7F821F6E475811E403E004FFBFE791FF061DE07FF3AF8C80F5D1B9EC1B6;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h0DC000157DEA07DB79A761FFEADDB0137FF8CC78B60FA0022FB19EABFEF05415;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h7F6939493BFC7FE596770069002844FF2041FFCC16EFFFCF91811BEFF181B460;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h78F170C0A1C29EBFFCD44BFD9D8E4A7403FACE03604F937FB7EF077F537B0939;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h2F3D8A1936043EB1D6F10F8C64C60FF783C7FFEA6B1DFFB8A218081AEFA58414;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h177FADC1FC755EFDFB4AA7FCBBE44B5118EFF75CBA77A57B64C3DCC61FF7A39C;
defparam sdpb_inst_1.INIT_RAM_22 = 256'hEFF8C014001F8FED1EF484B7EE903FC70044FF8243D7FE8C000C003C17ABFBC6;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h3D7684017C01C4DE81E707FD8743C401737F43ADE8ABD19900E040B370FE7C9A;
defparam sdpb_inst_1.INIT_RAM_24 = 256'hFF0BA6A487C3C9CFF769A60CF8201380095FFE02B3FBF4CD00441F65A63FFF90;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h69FF0043D20025803FE373BA787DFDFC645C5DFA69443FC0022F014321018770;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h6277EFFFFDC8687F3818587DFC0DAFFC03200146F95107B7BEBF2DC4D5FFD541;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h03FFEFEFFEF7BBC974ED0025BEFDF57B8D05A8B70AC7F6E2A97F759EC07AA2C0;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h04DFFF4B09390109D37C801FE9E83FBF6B90DFE393021F7FDE31A6D8180D9EF4;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h001FADCBFF70FFFF1AB4FEBF7E86D60C10001E2E7C056FE78B9CDEE8BFF1C8D8;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h57F5C18FC430203A73F94001AD7187DAA379102412E3FFC14D7A73800297D6B5;
defparam sdpb_inst_1.INIT_RAM_2B = 256'hE901C42C676B5528DD3991EFC99C640D504FA7D1C8D0887B36C405B5BC897AC6;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h771D70EBD0EFF012F0FEFFB7EE93E69D150007541B67EB7F2762CBCFFFD34F8D;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h3F8D7A178F0028DF9571BFD05D3589CFFF6E03C7FFFC07A447383100005DC6FB;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h00BE5D9C33FC38A7F590094F5E5F31782F77F07EB9EB5F7071627FF20700BF80;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h1E277F1826DBEDDEBC40839A1F28FE1E87D90C0017FF90534383C73F7FF6A31D;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h6CB792741017F74C801646AB30E8602ED51AF8850452C148C82400771AE050FF;
defparam sdpb_inst_1.INIT_RAM_31 = 256'hF037E8760FB4008204FC5FE5B2196805DD527314D4FAC110A143F2D00FA2AEBD;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h5047E87086D18D26FE276A25039D28680000010FAC6503511E00248AF71FFA97;
defparam sdpb_inst_1.INIT_RAM_33 = 256'hDFBF2502E2BBB81AE047C089F1A9DAD4F571FF0B967C76D5C8F80002880A0D8A;
defparam sdpb_inst_1.INIT_RAM_34 = 256'hB01C447E4F4FF8AC37E85E114E300EFDFD4AFA3C7E221E6CDBF38E5F2FF5A6BC;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h03B77FB6101765D142570C23C401EDB5098ECE409AF0B53F3A011EFFB702BBB9;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h6B67007BFEC6E00D04D6A8FC4E7C901491044DF9A2E3E5F0439F2BDC14CC6272;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h1F634688AC845F9D0BCAF9F85BEE6DC2CF83ED820D490FEB7AF9102A0794977A;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h427DE1BE20CF7F06617253647CE6C7FF27F591F07C13E37FE44BCCF8694A116A;
defparam sdpb_inst_1.INIT_RAM_39 = 256'hF8B95FAC9CDF7FEB2C8896C4E077969C836066A5D7639066DCBFFFFE006E8CB4;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h8017AD2587506BEC53A82484697091B3ED03D6AA920C1119F8F6C0401ED8BBBB;
defparam sdpb_inst_1.INIT_RAM_3B = 256'hC344866A089B67E946FD5CCDF6A84F5C79AF6F38A9535FB28105CC005BAF3467;
defparam sdpb_inst_1.INIT_RAM_3C = 256'hFFCFE0B0B5FF6B1A4A470042635E75356EDF32B0F76A7877DB43F3AFEB48EC76;
defparam sdpb_inst_1.INIT_RAM_3D = 256'hBFBE3D007E91B308809FEA40D8E473394640CB4DA4B7DE2F7BBDFD9BE06B78F7;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h279025E0580B86FCF1D6CA47210C89A158B33B65BC00AEE2DAC000000F2EAA97;
defparam sdpb_inst_1.INIT_RAM_3F = 256'hF0A5CF341CFDFFFC0C0FEB5E00E7CA07EC9FE5A80C7FAA3A4381826F4EE0EC11;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b1;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'h7FFD2C5077CFFFFF0603EE91B40007FFD0000000FFFFFFB73CFDBFFFFB04005A;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h000004FFFE000040000D7BFA10010119F7FFFBD417DCA08004DFFD0010000A7F;
defparam sdpb_inst_2.INIT_RAM_02 = 256'h0800000448FFFFFFF4F3C000008FFFC4032E00124E470000030607FFFFD660BF;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h00001FFF00417E34117F5000000028CDFFFFFFEA0E000023FFD401E1800003FA;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h000B20018F79FFFFFFC0100023FFFC081D817FD7EDA008000004FBFFFFFEE900;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h0003BFF858FCBC4DFFFF8000000007FBFFFFFFFE000001AFFFA083BC2FFFFED0;
defparam sdpb_inst_2.INIT_RAM_06 = 256'h4EE00602EFDFFDFFFE0000005FFB70CBBDAC7FFFF007D001801E37FFFFFFE800;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h05B7ECC0FBFDC71FFFD0190D10000FFDFFFFFFE0000047FFFC021F517BBFFD00;
defparam sdpb_inst_2.INIT_RAM_08 = 256'h7C600003AFFB5FFFE0000017FFFBBBF0FFBB01FD02960C00007BFDFFFFFE0001;
defparam sdpb_inst_2.INIT_RAM_09 = 256'h52DFF9AAE4FE80C0760377A9000046FFFFFFFE200003FFFFFF7DD7FE380F64BC;
defparam sdpb_inst_2.INIT_RAM_0A = 256'h90E0222EBFFE6DFE00805FFFFFCE6CE75D3F87C83C433804841EF7FEDFE00013;
defparam sdpb_inst_2.INIT_RAM_0B = 256'hFFFFE309FE01B8CFFFBC881E00005FEFFE9EE0004BB7FFFD375ED41A18FF69EF;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h2A80003B7F7DBFE00031FFFFF8A0DFFA0BEC7FF1EE65300008558C3BF600020F;
defparam sdpb_inst_2.INIT_RAM_0D = 256'h77F10861A26EFA1219E0E236000A1DFD6B7E0101528FFF474FD2422041C3CF42;
defparam sdpb_inst_2.INIT_RAM_0E = 256'hF7C00577F8B9BE0002200A3F1CA7C8228EC18AE94AEEB0000FBED55FE00A5839;
defparam sdpb_inst_2.INIT_RAM_0F = 256'h641587E3376183F5B01419D7602FFC40FFE000040253C3888E0E760C3DD374F9;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h71A2BFFFE06FE00100A8C3B1042866CD7853A7363578EE0BAEEF42BE00010042;
defparam sdpb_inst_2.INIT_RAM_11 = 256'h46B40007F2EFFC9FF025017EFFDF5B68FF80100960A1238156E759DEC8FC71BD;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h8067FF71E9FF80000A4442D6DB001F94FEE1FF41392C0EBEFEFB3AF000002B58;
defparam sdpb_inst_2.INIT_RAM_13 = 256'h49118B942CFC12FE111D20171FF69EB1F40000031FBA4F046991CFC94FF570B9;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h0987FD9E07F9100041FBA98FE02F749F2C2FA771F04311FFE5456F10000073F8;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h8FFA0B333C15295BC1750119FFB78D9FA000077FA56000046C93E3F5325C5890;
defparam sdpb_inst_2.INIT_RAM_16 = 256'hE53FFE6EFF80020FFA28E5C1B5ECC7C0BB58FDE6C00773FF9C57FA0024BF33C7;
defparam sdpb_inst_2.INIT_RAM_17 = 256'h7FFA7D1E003564DFE06928B3FFEFC7FE0003F8582D53824E18FC01F3813EF631;
defparam sdpb_inst_2.INIT_RAM_18 = 256'h33FF7C0EF80007F12A0C2680F007C001B243FF7445513FF9D23F90007F048E0C;
defparam sdpb_inst_2.INIT_RAM_19 = 256'hFFFFFF8007001FDF981E09BFFF147F80417E35BE3CC0FFEAE000038DFEFBAAC2;
defparam sdpb_inst_2.INIT_RAM_1A = 256'h9EFDD07FC000278ACAEA0FDFFEC00040DFFFBE2F4163F7CCDDFC008DF9DD8758;
defparam sdpb_inst_2.INIT_RAM_1B = 256'h23C8000053961DFFC603A4FBE88FF80044FC692661FCFFC400007F7C2DF35EEE;
defparam sdpb_inst_2.INIT_RAM_1C = 256'hF7E4E7D801F6FF8606B2C03E000004001BFFFF845ECFFF3AFFC80F5FE32E598E;
defparam sdpb_inst_2.INIT_RAM_1D = 256'h50C000110715FFFFFE83F3FFEADFB0177FFF0F85CE0FE000000121A7FFFF88C7;
defparam sdpb_inst_2.INIT_RAM_1E = 256'hFF693FE93BFC7FF9578F086B003CC000DFFFFFF5327FFFCFF9811BEFFE0974E0;
defparam sdpb_inst_2.INIT_RAM_1F = 256'h78FF108126AD3D7FFEFD2FFD9DFE4A7403FF1B76E00F937770000082AF7FD1EB;
defparam sdpb_inst_2.INIT_RAM_20 = 256'hEF3FFE0936043F36BDF1CF9EDCC7557737BFFFF030FFFFBFA218081AF248DC10;
defparam sdpb_inst_2.INIT_RAM_21 = 256'h67FFD2C006B2F13DFCF98FFEBDE44B5118F5063CBC73877BC3C023263FF7C663;
defparam sdpb_inst_2.INIT_RAM_22 = 256'hEFFFC014001FEDF8FEF48A97FDF000ECFF33FFFA223FFFFC000C043F7207FBA6;
defparam sdpb_inst_2.INIT_RAM_23 = 256'hFEBE800053FFF37FFF9B1FFDFF43C4017D285FEDFB0FDBF9001FBFFCC2FFC05F;
defparam sdpb_inst_2.INIT_RAM_24 = 256'hFFFBA6A487F0B0BFF7FD9FC3F820067FFF8DFFF7B67FFFCD00441FAC19FFFFF4;
defparam sdpb_inst_2.INIT_RAM_25 = 256'hDFFF00622DFFC97FC6BFCFFDF87DFDFF0E93FDFFF3F1FFC00260FFFC7FFEAF67;
defparam sdpb_inst_2.INIT_RAM_26 = 256'hFDF7EFFFF09527FFFED7A3FFFC0E0003FCEFFE8FA4FFFFB7BEBFC49E3FFFE73F;
defparam sdpb_inst_2.INIT_RAM_27 = 256'hFFFFEEF80108743685363FDDBFFFFE5DDCFFFFC2F53FFFE2AA008A66FF8439F7;
defparam sdpb_inst_2.INIT_RAM_28 = 256'hFFDFFFF585F0FFFE40917FFFE9FE8040904F204EBEFDFF7FFFDA9747FFF34093;
defparam sdpb_inst_2.INIT_RAM_29 = 256'hFFFFAA5400850000177E017F7FF8F7F2AFFFEA1293FFFFE74063214D4003B5F7;
defparam sdpb_inst_2.INIT_RAM_2A = 256'hFFFF18BC4E8FDFDE07A6BFFFFD533824808000B54D1FFFFE4DDF687FFCE0464A;
defparam sdpb_inst_2.INIT_RAM_2B = 256'h16FFF19036988008FAC70FFFF3170184AFB06094372F7FFA743B4B00000F8F69;
defparam sdpb_inst_2.INIT_RAM_2C = 256'hFFEB4F84141003C3D80100001039BA87040006F6C2FFFC63B88544303A1CC072;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h3E2A0B873F0028DF8A067FFCD9E914C0004428C0000007F436F9700000543327;
defparam sdpb_inst_2.INIT_RAM_2E = 256'hFB21E814700038D0F1000E97E05F0FF82F77F60147FF9CCE2F160004853C0000;
defparam sdpb_inst_2.INIT_RAM_2F = 256'hA0A81B07FEDBFFFF73CFFC8BC71C760000DDDC0007C5AFA5C07FC77FFFE01EFF;
defparam sdpb_inst_2.INIT_RAM_30 = 256'h6E02CFEC0019FA5C801791A3ADD81FEFFFFFFE1EFF8BD3EEB0E000F7DDE010F0;
defparam sdpb_inst_2.INIT_RAM_31 = 256'h80320D01FFFFFFFFFA0053A00F2CE005BEA5F314E61D23C2A0BFFFFFFFF24143;
defparam sdpb_inst_2.INIT_RAM_32 = 256'hFF77CBF086AE1CF6FFC99DC70E4407FFFFFFFFE0272716948E0033F0CF1FFCCE;
defparam sdpb_inst_2.INIT_RAM_33 = 256'hD9BFCE001D4447E5009251A99C9FDAFA074FFFF35F7077D78007FFFD77F40D7E;
defparam sdpb_inst_2.INIT_RAM_34 = 256'hB0633FFF950E47FFC6C1D6014EA2010202B50433C81A075BFBFDA016FFFE31AE;
defparam sdpb_inst_2.INIT_RAM_35 = 256'h84EFBAF60000000175C8DC0FB3FFF011D07FF06FFA8203CA8A00010040072881;
defparam sdpb_inst_2.INIT_RAM_36 = 256'h1AC0FF821F2E1FF169D542930F5FF00400005EE800006D0FFC0137C3FB0E8F1A;
defparam sdpb_inst_2.INIT_RAM_37 = 256'hDB7CB417EC805FFE7011077E041057F9C07C0EE72AB5D80879F9102007E38000;
defparam sdpb_inst_2.INIT_RAM_38 = 256'h2E0001C5DDC0000727E19E644D01FFFF27FFE4EF83B4A00007FDFC07816B72E5;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h70D045B3FFFFFFD2ACD5A740007ECB8C00007597F71D1EDB147FFFFFFF523EA2;
defparam sdpb_inst_2.INIT_RAM_3A = 256'h8017C5A2DF506BF137D6128546810FEFFFFC1D2E8CBC011EF059C0001F33D1BD;
defparam sdpb_inst_2.INIT_RAM_3B = 256'h05C9A1A5F7641A0A6D793CCDF84B5CFC79AF8A45C88B3CD494FF7FEFA4C2D0F5;
defparam sdpb_inst_2.INIT_RAM_3C = 256'hFFF2762DFFFFFFE3E692F7E4B95C0A4A91213CC38F6AFFB2275BF3AFFC69CF52;
defparam sdpb_inst_2.INIT_RAM_3D = 256'h8D87CB8000001109FFFFFFFF16E35FFFFFFF0D90169C84A1D0000000007007F7;
defparam sdpb_inst_2.INIT_RAM_3E = 256'hD840329FA7F47900E51941F65E4C088040B33FFFFFFF50E201FFFFFFF0330F57;
defparam sdpb_inst_2.INIT_RAM_3F = 256'h4A7E5F341CFFFFFFFFF0048000A035F8136001D0369BD7C4C101026F4EFFFFEE;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b1;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'h7FFD2C5077CFFFFFFFFC016E4BFFFFFFD0000000FFFFFFB73CFDBFFFFFFFFFA2;
defparam sdpb_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFE000FC0000D7BFA10010119F7FFFFFFE8235F7FFFFFFD00F0000A7F;
defparam sdpb_inst_3.INIT_RAM_02 = 256'h0800000448FFFFFFFFFC3FFFFFFFFFC007FC00124E470000030607FFFFFFFF40;
defparam sdpb_inst_3.INIT_RAM_03 = 256'hFFFFFFFF007EAFE4117F5000000028CDFFFFFFFFF1FFFFFFFFD4012F5C0003FA;
defparam sdpb_inst_3.INIT_RAM_04 = 256'h000B20018F79FFFFFFFFEFFFFFFFFC0FFDFF7FD7EDA008000004FBFFFFFFFEFF;
defparam sdpb_inst_3.INIT_RAM_05 = 256'hFFFFFFF835CF6CFFFFFF8000000007FBFFFFFFFFFFFFFFFFFFA0FEDFF6FFFED0;
defparam sdpb_inst_3.INIT_RAM_06 = 256'h46200602EFDFFDFFFFFFFFFFFFFB7FDDFFFFEFFFF007E001801E37FFFFFFF7FF;
defparam sdpb_inst_3.INIT_RAM_07 = 256'hFFFFFCBFC9F3CFFFFFD0117D10000FFDFFFFFFFFFFFFFFFFFDFFDFCEFFFFFD00;
defparam sdpb_inst_3.INIT_RAM_08 = 256'h83E00003AFFB5FFFFFFFFFFFFFF871E47F87FFFD03297400007BFDFFFFFFFFFE;
defparam sdpb_inst_3.INIT_RAM_09 = 256'hFFFFFB9FEBFF3F3FF603F82B000046FFFFFFFFDFFFFFFFFFF27F9FF8F7FF64BC;
defparam sdpb_inst_3.INIT_RAM_0A = 256'hEFE0222EBFFE6DFFFFFFFFFFFFD87DE37BD07FC83BB8D804841EF7FEDFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0B = 256'hFFFFE7F9FF1E783FFFBECA7E00005FEFFE9EFFFFFFFFFFFFFD6ECFFD07FF69CA;
defparam sdpb_inst_3.INIT_RAM_0C = 256'hF780003B7F7DBFFFFFFFFFFFFFEF0FD5FFE3FFFFF752F00008558C3BF7FFFFFF;
defparam sdpb_inst_3.INIT_RAM_0D = 256'hFFFE75DD5E2F35FD7DBE3FFE000A1DFD6B7FFFFFFFFFFFFE3D91BCEE3FFB0F83;
defparam sdpb_inst_3.INIT_RAM_0E = 256'hFBC00577F8B9BFFFFFFFFFFFE7EA2F9FEA3E19AC72FFB0000FBED55FFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0F = 256'h3EE2FF1E7E687DF044E9FBAF602FFC40FFFFFFFFFFFFFC57D17DEE43CFED3005;
defparam sdpb_inst_3.INIT_RAM_10 = 256'h89AABFFFE06FFFFFFF59E7AE79D7CDECC7871FD3CE5C9E0BAEEF42BFFFFFFF7E;
defparam sdpb_inst_3.INIT_RAM_11 = 256'hF8DBDF7FEA60267FF84B3BB1FFDF5B68FE7FFFFD8F79C20E8FDFD4222FFF7C77;
defparam sdpb_inst_3.INIT_RAM_12 = 256'h7F9FFF71E9FE7FFFFD41411B15F39F0C03F7FFA6C87BF3BEFEFB3AEFFFFF8463;
defparam sdpb_inst_3.INIT_RAM_13 = 256'h71F746CF1C01E1FF85EEDFE8FFF69EB1EBFFFFF01F8392F76EB0C0003FFA9E62;
defparam sdpb_inst_3.INIT_RAM_14 = 256'hF67FFD9E07E6EFFFBE252E0FCFBE7380C99FF0EEC5BCEBFFE5456EEFFFFF839A;
defparam sdpb_inst_3.INIT_RAM_15 = 256'h80039B0F03E2266E7E7EFEE4FFB78D9E5FFFF88D808000B9EC701C88FC39EC6F;
defparam sdpb_inst_3.INIT_RAM_16 = 256'h16FFFE6EFE7FFDF006CD9C3E36E3C03F22C77BF3BFF8EFFF9C57E5FFDB40E4E7;
defparam sdpb_inst_3.INIT_RAM_17 = 256'hFFF87D01FFD35CBFFBC3D7AFFFEFC7E1FFFC00A41CCFFC21F803FB240EFF75EE;
defparam sdpb_inst_3.INIT_RAM_18 = 256'hEFFF7C0EE7FFF801AC469E8000003FFE1C9FFFACD44EFFF9D23E6FFF80095125;
defparam sdpb_inst_3.INIT_RAM_19 = 256'h0000007FFFFFFFDFECFA7B7FFF147E7FBE8038002BC000001FFFFC0BFEFD46E3;
defparam sdpb_inst_3.INIT_RAM_1A = 256'hFEFDD07E3FFFD80C9BA60020013FFFFFFFFFBFB54F67F7CCDDE3FF7201945D38;
defparam sdpb_inst_3.INIT_RAM_1B = 256'hDC37FFFFFFFF67FFF84375FBE88FE7FFBB00739DE003003BFFFFFFFFEDFC68FB;
defparam sdpb_inst_3.INIT_RAM_1C = 256'hF7E4E7E7FE090007FFCE3FC1FFFFFFFF90BFFFF81DFFFF3AFE37F0A003CE3981;
defparam sdpb_inst_3.INIT_RAM_1D = 256'hBFBFFFE7F4FFFFFFFF53F3FFEADE4FE880000FF2A1F01FFFFFFE725FFFFFE2C6;
defparam sdpb_inst_3.INIT_RAM_1E = 256'hFF693E16C403800188E0F796FFC53FFFFFFFFFFAAFDFFFCFE67EE410000EAA1F;
defparam sdpb_inst_3.INIT_RAM_1F = 256'h87020F7E7990217FFFBC7FFD9DE1B58BFC0011DA1F706C878FFFFFFCE77FF5BF;
defparam sdpb_inst_3.INIT_RAM_20 = 256'hEF3FE1F6C9FBC02B5C0E704073389F0825C7FFFB39FFFFBE5DE7F7E50322C3E7;
defparam sdpb_inst_3.INIT_RAM_21 = 256'h0700023FF853283DFEB37FFEBE1BB4AEE7063F0343883484643FD7EE8FF7DDFF;
defparam sdpb_inst_3.INIT_RAM_22 = 256'hEFFE3FEBFFE00AAC010B40480B8FFF13FFE2FFF5EC7FFFE3FFF3FBC071A00439;
defparam sdpb_inst_3.INIT_RAM_23 = 256'h00117FFE0FFFFBBFFD50FFFDE0BC3BFE81CBC012184822C6FFE07FFECAFFBB23;
defparam sdpb_inst_3.INIT_RAM_24 = 256'hFFE4595B7803E5800800C02007DFE7FFFFE9FFE0A9FFFE32FFBBE0368800001A;
defparam sdpb_inst_3.INIT_RAM_25 = 256'h4000FF95FFFFF0FFF8603FFE0782020051F002007800003FFC1FFFFE1FFF1187;
defparam sdpb_inst_3.INIT_RAM_26 = 256'hFE081000014360000050200003F09FFFFF27FFF1C3FFE04841400B4200000601;
defparam sdpb_inst_3.INIT_RAM_27 = 256'h00001037FFFF93FFFC08FFE2400000665400001E0680001D49FFFFFC7FFF832F;
defparam sdpb_inst_3.INIT_RAM_28 = 256'hE02000062CE8000058110000160E7FFFFEFFFF8251FE0080001C90C0000240E0;
defparam sdpb_inst_3.INIT_RAM_29 = 256'h000051DFFFF8BFFFE4117E008001A85580000C033000001833FFFFA7FFFC880F;
defparam sdpb_inst_3.INIT_RAM_2A = 256'h000018BCE580001C06E000000287FFFF5FFFFF6423E000004DA2580000907A00;
defparam sdpb_inst_3.INIT_RAM_2B = 256'h0000046FCA97FFF70822E000031E41DC0001E0EC00000004B3FFA1FFFFF1143E;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h000F67A09C0002C32800000000315FBEFBFFF8444C0000433B0EC0002E18C000;
defparam sdpb_inst_3.INIT_RAM_2D = 256'h3FCBCBD680FFD72010400000DDED0F40004C3DC0000007E0D4040FFFFFA00040;
defparam sdpb_inst_3.INIT_RAM_2E = 256'h028DC47EF00068EBF1000FE47FDF0007D08809A0200013FC805E000686DC0000;
defparam sdpb_inst_3.INIT_RAM_2F = 256'h2855DB0001240000600000D3CF840E0001DFBC0007F909F8C0003880000C0200;
defparam sdpb_inst_3.INIT_RAM_30 = 256'hBE063BDC001FFCBC8017E41C46A80010000003A4001A0329A9E00097EBE010FF;
defparam sdpb_inst_3.INIT_RAM_31 = 256'h7FC8D700000000000000AF63017BE0051FDBF314F8B3DF1B2000000000020001;
defparam sdpb_inst_3.INIT_RAM_32 = 256'hCE64C7F0875FDBF6FFF2EF9CD06C0000000000002933262F7E0031FDBF1FFF13;
defparam sdpb_inst_3.INIT_RAM_33 = 256'hAE5078000000000000F21109A27FDAE5FA3FFFFC7D7B80B18000000000000F0E;
defparam sdpb_inst_3.INIT_RAM_34 = 256'h305EFFFFE0F53FFFF8B9F1FEB1DE000000000039C4160CA7FBFE9FA1FFFFC476;
defparam sdpb_inst_3.INIT_RAM_35 = 256'h7FF7C7EE000000017DC00002EFFFFECE77FFFF89FA1FFBF20A0000000007B800;
defparam sdpb_inst_3.INIT_RAM_36 = 256'h029FFFFD4001FFFE898693610FB4700400005F38000014FFFFE4C73FFFF09136;
defparam sdpb_inst_3.INIT_RAM_37 = 256'h0080D5EFEC805FFFA8000085FFFF840A3FFFF0841606200CCFF9102007FB8000;
defparam sdpb_inst_3.INIT_RAM_38 = 256'hC9FFFE34103FFFF85827369B8A127FFF27FFF92000511FFFF941E3FFFE8F8D9E;
defparam sdpb_inst_3.INIT_RAM_39 = 256'hAF14D0AFFFFFFFFCC8CBF33FFF8543C3FFFF86572F42E0C0B7FFFFFFFF95115A;
defparam sdpb_inst_3.INIT_RAM_3A = 256'h7FE80CE7C0AF9401AAB34479DF51FFFFFFFFE69E56A3FEE0EC6C3FFFE02799FC;
defparam sdpb_inst_3.INIT_RAM_3B = 256'h467E11BFFFFFFFF4766B0332009FCC0386500C81EEC0BDE497FFFFEFFF0AB9BC;
defparam sdpb_inst_3.INIT_RAM_3C = 256'h00033F74000000038F57745DD817FFFFFFFEC0FF8095003277440C500073CFFE;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h44520F7FFFFFEEF60000000019F6C00000000E3F928949812FFFFFFFFF800008;
defparam sdpb_inst_3.INIT_RAM_3E = 256'h0000318000000000F8E1476A0063F77FBF4CC000000000E378000000003C925F;
defparam sdpb_inst_3.INIT_RAM_3F = 256'hF80050CBE30000000000000000E00000000001E7C5F518063EFEFD90B1000000;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b1;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'h7FFD2C5077CFFFFFFFFFFFFFFFFFFFFFD0000000FFFFFFB73CFDBFFFFFFFFFFE;
defparam sdpb_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFE000FC0000D7BFA10010119F7FFFFFFFFFFFFFFFFFFFD00F0000A7F;
defparam sdpb_inst_4.INIT_RAM_02 = 256'h0800000448FFFFFFFFFFFFFFFFFFFFC003FE00124E470000030607FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_03 = 256'hFFFFFFFF005DB7E4117F5000000028CDFFFFFFFFFFFFFFFFFFD401EFD80003FA;
defparam sdpb_inst_4.INIT_RAM_04 = 256'h000B20018F79FFFFFFFFFFFFFFFFFC07FAFF3FD7EDA008000004FBFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_05 = 256'hFFFFFFF87DFFAFFFFFFF8000000007FBFFFFFFFFFFFFFFFFFFA1FEABF7FFFED0;
defparam sdpb_inst_4.INIT_RAM_06 = 256'h56600602EFDFFDFFFFFFFFFFFFFB7FBDFCBFDFFFF007B001801E37FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_07 = 256'hFFFFFCDFEFF5DAFFFFD01FBB10000FFDFFFFFFFFFFFFFFFFFDFF5FD3FDFFFD00;
defparam sdpb_inst_4.INIT_RAM_08 = 256'h3FA00003AFFB5FFFFFFFFFFFFFF97DFCBFFFFFFD037A7400007BFDFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_09 = 256'hFFFFFB9FED7EAEFFF603AFFB000046FFFFFFFFFFFFFFFFFFB57FE7FFFFFF64B6;
defparam sdpb_inst_4.INIT_RAM_0A = 256'h91E0222EBFFE6DFFFFFFFFFFFFDFFD654EEFFFC83CFA1804841EF7FEDFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0B = 256'hFFFFFEF7FEBEF7FFFFBFE00600005FEFFE9EFFFFFFFFFFFFDF2ED7E9FFFF69EC;
defparam sdpb_inst_4.INIT_RAM_0C = 256'h6180003B7F7DBFFFFFFFFFFFFE9F7FFDCF1FFFFFFA04300008558C3BF7FFFFFF;
defparam sdpb_inst_4.INIT_RAM_0D = 256'hFFFF73FF7CEF0FFE76FF600E000A1DFD6B7FFFFFFFFFFFFF7E5D9AE1FFFF8BE8;
defparam sdpb_inst_4.INIT_RAM_0E = 256'h01C00577F8B9BFFFFFFFFFFFFF23E78EE9FFF57EFA0070000FBED55FFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0F = 256'hFFFA3E7EDF67FEF3F97E043F602FFC40FFFFFFFFFDFFFFF3BFFBE63FF721DEC2;
defparam sdpb_inst_4.INIT_RAM_10 = 256'h09AABFFFE06FFFFFFFBFEF5FBDFBDDED3FEE7FE2F0A1FE0BAEEF42BFFFFFFF7D;
defparam sdpb_inst_4.INIT_RAM_11 = 256'h1F0DBF7CF21FDAFFFCFC83DFDFDF5B68FFFFFFFEDFFFFF8DCBE653FCB7FFC981;
defparam sdpb_inst_4.INIT_RAM_12 = 256'hFFFFFF71E9FFFFFFFFBFBFE3FEF7BE03FDFFFFC9E4F7FFBEFEFB3AFFFFFFFFAC;
defparam sdpb_inst_4.INIT_RAM_13 = 256'h81F7D5CF03FE37FFDCF6FFFFFFF69EB1FFFFFFF7E07C1EEF24B03FEEFFFCAF1B;
defparam sdpb_inst_4.INIT_RAM_14 = 256'hFFDFFD9E07FFFFFFFF88C00FCF9F707FFBBFF9BF5DFFFBFFE5456FFFFFFFFC1B;
defparam sdpb_inst_4.INIT_RAM_15 = 256'h8003BF00FFFA9FB9BFFFFFFFFFB78D9FFFFFFFFF3F80003FEC0FFF73FF5FF4FF;
defparam sdpb_inst_4.INIT_RAM_16 = 256'hF5FFFE6EFFFFFFFFFE2F7C003FE03FFFFDAEE7F9FFFFFFFF9C57FFFFFFFFF4F7;
defparam sdpb_inst_4.INIT_RAM_17 = 256'h000782FFFFE5747FFDBFFF9FFFEFC7FFFFFFFFE7F3C0001007FFFC3375FFBBFF;
defparam sdpb_inst_4.INIT_RAM_18 = 256'h1FFF7C0EFFFFFFFE4F9D817FFFFFFFFFDFFFFFCFFDBDFFF9D23FFFFFFFF47E9C;
defparam sdpb_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFDFF1A705FFFF147FFFFFFFC1FF983FFFFFFFFFFFF7FEFE46FC;
defparam sdpb_inst_4.INIT_RAM_1A = 256'h7EFDD07FFFFFFFF0F761FFFFFFFFFFFFFFFFBFC6201FF7CCDDFFFFFFFE190B07;
defparam sdpb_inst_4.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFF9401FBE88FFFFFFFFF827C1FFFFFFFFFFFFFFFEDFF8C42;
defparam sdpb_inst_4.INIT_RAM_1C = 256'h77E4E7FFFFFFFFF80041FFFFFFFFFFFFC37FFFFEA10FFF3AFFFFFFFFFC0E067F;
defparam sdpb_inst_4.INIT_RAM_1D = 256'hFF7FFFF803FFFFFFFFA82FFFEADFFFFFFFFFF01D1FFFFFFFFFFFCDFFFFFFF531;
defparam sdpb_inst_4.INIT_RAM_1E = 256'hFF693FFFFFFFFFFE525FFFFFFFF3FFFFFFFFFFFD703FFFCFFFFFFFFFFFF085FF;
defparam sdpb_inst_4.INIT_RAM_1F = 256'hFFFE3FFF9EDF7AFFFF439FFD9DFFFFFFFFFFE7B1FFFFEFF97FFFFFFF3F7FEA61;
defparam sdpb_inst_4.INIT_RAM_20 = 256'hEF3FFFFFFFFFFFC3D3FFFFDF6FFF44FFF7FFFFFE847FFFBFFFFFFFFFFC6EBFFF;
defparam sdpb_inst_4.INIT_RAM_21 = 256'hF2FFF9FFFC6C783DFF8A1FFEBFFFFFFFFFF8B2FFFBFBC3FFABFFF7EE0FF7F313;
defparam sdpb_inst_4.INIT_RAM_22 = 256'hEFFFFFFFFFFFF3EBFFFDDFBFF57FFF87FFB3FFFC19FFFFFFFFFFFFFFA21FFFFF;
defparam sdpb_inst_4.INIT_RAM_23 = 256'hFFEFFFFF1FFFFB3FFF011FFDFFFFFFFFFE573FFFE7A7FFBFFFF0FFFFCAFFE063;
defparam sdpb_inst_4.INIT_RAM_24 = 256'hFFFFFFFFFFFCF07FFFFE3FD7FFFFF3FFFFF9FFF081FFFFFFFFFFFFC7E7FFFFE5;
defparam sdpb_inst_4.INIT_RAM_25 = 256'hFFFFFFE1FFFFF4FFFC463FFFFFFFFFFFABCFFFFF87FFFFFFFF1FFFFF1FFF810F;
defparam sdpb_inst_4.INIT_RAM_26 = 256'hFFFFFFFFFE141FFFFF0FDFFFFFFE9FFFFFEFFFE1C9FFFFFFFFFFF159FFFFF8FE;
defparam sdpb_inst_4.INIT_RAM_27 = 256'hFFFFFF7FFFFFF7FFF8087FFFFFFFFF86D3FFFFE5FA7FFFFFF8FFFFFA3FFF000F;
defparam sdpb_inst_4.INIT_RAM_28 = 256'hFFFFFFF81927FFFFA7E4FFFFFFF6FFFFFC3FFFE603FFFFFFFFE0963FFFFCBF2F;
defparam sdpb_inst_4.INIT_RAM_29 = 256'hFFFFFDDFFFFC7FFFFC00FFFFFFFEFE747FFFF2FCCFFFFFFF93FFFFC3FFFF861F;
defparam sdpb_inst_4.INIT_RAM_2A = 256'hFFFFE8B90C7FFFEDFB9FFFFFFFEFFFFF87FFFFE407FFFFFFCD75C7FFFF2F81FF;
defparam sdpb_inst_4.INIT_RAM_2B = 256'hFFFFFBEFF28FFFFFF803FFFFFD1C1143FFFE5F33FFFFFFFF17FFF17FFFFF111F;
defparam sdpb_inst_4.INIT_RAM_2C = 256'hFFF37F00F3FFFCBC67FFFFFFFFD6FFBDFFFFFFD44FFFFFA3EB0A3FFFD9E23FFF;
defparam sdpb_inst_4.INIT_RAM_2D = 256'hC00C04167FFFFFFFF003FFFF1FEB093FFF83C43FFFFFF8636BFCFFFFFFFC223F;
defparam sdpb_inst_4.INIT_RAM_2E = 256'hFCEFD41C0FFF87000EFFF0058060FFFFFFFFFFA81FFFE7ECE091FFF978C3FFFF;
defparam sdpb_inst_4.INIT_RAM_2F = 256'h37FE14FFFFFFFFFFE03FFF0FF68161FFFA2183FFF801D6023FFFFFFFFFFC01FF;
defparam sdpb_inst_4.INIT_RAM_30 = 256'h22060443FFE200837FE8062FB0D7FFFFFFFFFC43FFEC03E8541FFF48181FEF00;
defparam sdpb_inst_4.INIT_RAM_31 = 256'h7FD7B8FFFFFFFFFFFFFF6F6000881FFA00180CEB00FDFCC25FFFFFFFFFFDFFFF;
defparam sdpb_inst_4.INIT_RAM_32 = 256'hDF67E00F78C00809000337FBCDB3FFFFFFFFFFFFCFBF263101FFC40180E0001B;
defparam sdpb_inst_4.INIT_RAM_33 = 256'hF7ED9BFFFFFFFFFFFF3E8149B2002500010000006DFFFFE3FFFFFFFFFFFFF0EE;
defparam sdpb_inst_4.INIT_RAM_34 = 256'hB0F200000407000000DFFEEFFE71FFFFFFFFFFC3FC0E0F200400C0300000067E;
defparam sdpb_inst_4.INIT_RAM_35 = 256'hFB7FFD51FFFFFFFE81C02C05200000407000000DFAFDDFFCB5FFFFFFFFF83980;
defparam sdpb_inst_4.INIT_RAM_36 = 256'h03C00001C06000000CC181F10FD20FFBFFFFA07800401800000C01000000CB32;
defparam sdpb_inst_4.INIT_RAM_37 = 256'h2200FB40137FA0001800016400000C0E000000D74142000DF806EFDFF8018000;
defparam sdpb_inst_4.INIT_RAM_38 = 256'hF800003C1C0000006A3B9EC00E1D0000D80000E0003F800000C1A000000D5A03;
defparam sdpb_inst_4.INIT_RAM_39 = 256'h001FDB5000000000C43A5D000007C2C00000075FF0A800FF4A000000001B7805;
defparam sdpb_inst_4.INIT_RAM_3A = 256'h00000F6440000001C8F0F681BFFE80000000075E3EE0000084740000003AA9C3;
defparam sdpb_inst_4.INIT_RAM_3B = 256'hB73FFE40000000007867000000F7B40000000F2FF30C3BFA64000010000C612C;
defparam sdpb_inst_4.INIT_RAM_3C = 256'h0003EF9C00000003F5F78963E7AC0000000000FF80000034FCC00000007D67D1;
defparam sdpb_inst_4.INIT_RAM_3D = 256'hB3FDF30000000000000000001FFAC00000000FD791763F5E2000000000000000;
defparam sdpb_inst_4.INIT_RAM_3E = 256'h0000398000000000FEE17C9DBF80000000000000000000E328000000003F3A58;
defparam sdpb_inst_4.INIT_RAM_3F = 256'h03FFB000000000000000000000E00000000001FB8524C7F80000000000000000;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b1;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'h7FFD2C5077CFFFFFFFFFFFFFFFFFFFFFD0000000FFFFFFB73CFDBFFFFFFFFFFE;
defparam sdpb_inst_5.INIT_RAM_01 = 256'hFFFFFFFFFE001040000D7BFA10010119F7FFFFFFFFFFFFFFFFFFFD0090000A7F;
defparam sdpb_inst_5.INIT_RAM_02 = 256'h0800000448FFFFFFFFFFFFFFFFFFFFC0040200124E470000030607FFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_03 = 256'hFFFFFFFF0061D814117F5000000028CDFFFFFFFFFFFFFFFFFFD40170E40003FA;
defparam sdpb_inst_5.INIT_RAM_04 = 256'h000B20018F79FFFFFFFFFFFFFFFFFC080F00FFD7EDA008000004FBFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_05 = 256'hFFFFFFF84E30F303FFFF8000000007FBFFFFFFFFFFFFFFFFFFA101DC18FFFED0;
defparam sdpb_inst_5.INIT_RAM_06 = 256'h62600602EFDFFDFFFFFFFFFFFFFB707603C03FFFF007F001801E37FFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_07 = 256'hFFFFFCE0770E3D8FFFD0110310000FFDFFFFFFFFFFFFFFFFFE01E03F06FFFD00;
defparam sdpb_inst_5.INIT_RAM_08 = 256'h00600003AFFB5FFFFFFFFFFFFFFB8C1FC078FFFD03A00C00007BFDFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_09 = 256'hFFFFFBB017C181FFF603D01F000046FFFFFFFFFFFFFFFFFFBF8078040FFF64B9;
defparam sdpb_inst_5.INIT_RAM_0A = 256'h80E0222EBFFE6DFFFFFFFFFFFFDCC39FB02FFFC83F081804841EF7FEDFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0B = 256'hFFFFF6EE00A00FFFFFBF008600005FEFFE9EFFFFFFFFFFFFDFB13C00FFFF69FA;
defparam sdpb_inst_5.INIT_RAM_0C = 256'h6180003B7F7DBFFFFFFFFFFFFE8FB02620FFFFFFFD04300008558C3BF7FFFFFF;
defparam sdpb_inst_5.INIT_RAM_0D = 256'hFFFF71BF8102FFFF800FE20E000A1DFD6B7FFFFFFFFFFFFE7BEE001FFFFCF7F8;
defparam sdpb_inst_5.INIT_RAM_0E = 256'h83C00577F8B9BFFFFFFFFFFFFF33F84057FFE3911E1070000FBED55FFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0F = 256'hFEFA3D60021FFF07FE17042F602FFC40FFFFFFFFFBFFFFD3FE0001FFF8DE61E0;
defparam sdpb_inst_5.INIT_RAM_10 = 256'h064ABFFFE06FFFFFFFFFEFFFF9D71072FFF1FFFC38217E0BAEEF42BFFFFFFF7F;
defparam sdpb_inst_5.INIT_RAM_11 = 256'h7FEDCF8215FFE1FFFF1E00203FDF5B68FFFFFFFEFFFEFF95F030EFFF4FFFB5C1;
defparam sdpb_inst_5.INIT_RAM_12 = 256'h0007FF71E9FFFFFFFFFFFFFC7FF810FFFE8FFFE1F08800BEFEFB3AFFFFFFFFDE;
defparam sdpb_inst_5.INIT_RAM_13 = 256'hFE0B6028FFFF47FFE3FB00007FF69EB1FFFFFFFFFFFFE0F3124FFFF1FFFE5F84;
defparam sdpb_inst_5.INIT_RAM_14 = 256'h001FFD9E07FFFFFFFFFE0FF027C18FFFF47FFE1F920007FFE5456FFFFFFFFFE5;
defparam sdpb_inst_5.INIT_RAM_15 = 256'h7FFD80FFFFFF7FC07FB00003FFB78D9FFFFFFFF0C07FFFBE33FFFF8FFFA3F800;
defparam sdpb_inst_5.INIT_RAM_16 = 256'h0FFFFE6EFFFFFFFFF9D083FFC51FFFFFD0704FFC00001FFF9C57FFFFFFFF0B00;
defparam sdpb_inst_5.INIT_RAM_17 = 256'hFFFFFFFFFFFAD9FFFE8000FFFFEFC7FFFFFFFF98003FFFFFFFFFFE480BFFD000;
defparam sdpb_inst_5.INIT_RAM_18 = 256'h1FFF7C0EFFFFFFFFF06C7FFFFFFFFFFFE0BFFFF40203FFF9D23FFFFFFFFF8183;
defparam sdpb_inst_5.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFDFFEC802FFFF147FFFFFFFFEBF87FFFFFFFFFFFFFFFEFF9902;
defparam sdpb_inst_5.INIT_RAM_1A = 256'h7EFDD07FFFFFFFFF1D1FFFFFFFFFFFFFFFFFBFF8108FF7CCDDFFFFFFFFE158FF;
defparam sdpb_inst_5.INIT_RAM_1B = 256'hFFFFFFFFFFFF83FFFFF081FBE88FFFFFFFFFFC03FFFFFFFFFFFFFFFFEDFFF242;
defparam sdpb_inst_5.INIT_RAM_1C = 256'h77E4E7FFFFFFFFFFFFBFFFFFFFFFFFFFCCFFFFFF870FFF3AFFFFFFFFFFF1FFFF;
defparam sdpb_inst_5.INIT_RAM_1D = 256'hFF7FFFFC2FFFFFFFFFE463FFEADFFFFFFFFFFFF87FFFFFFFFFFFCBFFFFFFFC19;
defparam sdpb_inst_5.INIT_RAM_1E = 256'hFF693FFFFFFFFFFFBFBFFFFFFFF0FFFFFFFFFFFF311FFFCFFFFFFFFFFFFFABFF;
defparam sdpb_inst_5.INIT_RAM_1F = 256'hFEFC7FFFC2E0E5FFFFC097FD9DFFFFFFFFFFFEC7FFFFFFF9FFFFFFFF9F7FF840;
defparam sdpb_inst_5.INIT_RAM_20 = 256'hEF3FFFFFFFFFFFFD0FFFFFDF5FFFB3FF8807FFFE043FFFBFFFFFFFFFFF8A7FFF;
defparam sdpb_inst_5.INIT_RAM_21 = 256'hF1FFF3FFFF9F87FDFF880FFEBFFFFFFFFFFFE9FFFBFBCFFFC7FFE811FFF7F201;
defparam sdpb_inst_5.INIT_RAM_22 = 256'hEFFFFFFFFFFFFC07FFFFDF7FF8FFFFFFFFCDFFFC097FFFFFFFFFFFFFDD7FFFFF;
defparam sdpb_inst_5.INIT_RAM_23 = 256'hFF9FFFFFFFFFFCFFFF003FFDFFFFFFFFFFBEFFFFFF9FFCFFFFFFFFFF3AFFE063;
defparam sdpb_inst_5.INIT_RAM_24 = 256'hFFFFFFFFFFFE8BFFFFFE7FEFFFFFFDFFFFE7FFF0A0FFFFFFFFFFFFF95FFFFFF3;
defparam sdpb_inst_5.INIT_RAM_25 = 256'h3FFFFFFFFFFFFBFFFC663FFFFFFFFFFFD4BFFFFFCFF9FFFFFFFFFFFFFFFF8097;
defparam sdpb_inst_5.INIT_RAM_26 = 256'hFFFFFFFFFFE2FFFFFFFFE7FFFFFF7FFFFF9FFFE0C9FFFFFFFFFFFEF7FFFFF9FF;
defparam sdpb_inst_5.INIT_RAM_27 = 256'hFFFFFF8FFFFFCFFFF8007FFFFFFFFFF10FFFFFF3FCFFFFFFF7FFFFFDFFFF012F;
defparam sdpb_inst_5.INIT_RAM_28 = 256'hFFFFFFFFD49FFFFFEFFFFFFFFFF9FFFFFFFFFFC413FFFFFFFFFF65FFFFFE7FBF;
defparam sdpb_inst_5.INIT_RAM_29 = 256'hFFFFFE3FFFFFFFFFF400FFFFFFFE04C3FFFFFDFF3FFFFFFFCFFFFFFFFFFE8A9F;
defparam sdpb_inst_5.INIT_RAM_2A = 256'hFFFFF75763FFFFF7FD7FFFFFFFF0FFFFFFFFFFAC27FFFFFFB2993FFFFF9FF7FF;
defparam sdpb_inst_5.INIT_RAM_2B = 256'hFFFFFC13FD7FFFFFE802FFFFFEE1BF3FFFFF3FCFFFFFFFFF8FFFFEFFFFFD043F;
defparam sdpb_inst_5.INIT_RAM_2C = 256'hFFFC98DF4FFFFE7F9FFFFFFFFFE00043FFFFFF440FFFFFDCD6F1FFFFEFF9FFFF;
defparam sdpb_inst_5.INIT_RAM_2D = 256'hFFFFFFE9FFFFFFFFD003FFFFA316F4FFFFFFF3FFFFFFFFBF8003FFFFFFF8083F;
defparam sdpb_inst_5.INIT_RAM_2E = 256'hFF5337E1FFFFDFF7FFFFFFFBFFBFFFFFFFFFFE883FFFFA337F4FFFFCFF3FFFFF;
defparam sdpb_inst_5.INIT_RAM_2F = 256'hCFEBEFFFFFFFFFFFA03FFFEC1FFFDFFFFDFE7FFFFFFE5FFFFFFFFFFFFFF403FF;
defparam sdpb_inst_5.INIT_RAM_30 = 256'h15F9F33FFFF9FF7FFFFFF9FF372FFFFFFFFFFE0FFFF03C77ABFFFF9FE7FFFFFF;
defparam sdpb_inst_5.INIT_RAM_31 = 256'hFE0BCFFFFFFFFFFFFFFF909FFE27FFFFBFE7FFFFFF27F2DFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_5.INIT_RAM_32 = 256'h00D85FFFFF7FF7FFFFFC7FC03E7FFFFFFFFFFFFFF058D9C4FFFFFBFE7FFFFFE0;
defparam sdpb_inst_5.INIT_RAM_33 = 256'h8003E3FFFFFFFFFFFFE13E9649FFFFFBFCFFFFFF86FC007F5FFFFFFFFFFFFE01;
defparam sdpb_inst_5.INIT_RAM_34 = 256'hCF09FFFFF3F8FFFFFF0FE0003FD7FFFFFFFFFFFC243DF09FFFFFBFCFFFFFF8FA;
defparam sdpb_inst_5.INIT_RAM_35 = 256'h807FFCBFFFFFFFFFFE3FE1F89FFFFF3FAFFFFFF0FBC003FE7FFFFFFFFFFF8600;
defparam sdpb_inst_5.INIT_RAM_36 = 256'hFCBFFFFF3F9FFFFFF13790010FEBFFFFFFFFFF87FFFFCBFFFFFBFCFFFFFF1736;
defparam sdpb_inst_5.INIT_RAM_37 = 256'h2200C0BFFFFFFFFFC7FFFF93FFFFE3F5FFFFFF18FF49000E0FFFFFFFFFFE7FFF;
defparam sdpb_inst_5.INIT_RAM_38 = 256'h67FFFFD3E3FFFFFF8CDFFEC00DE1BFFFFFFFFE1FFFF17FFFFE3E1FFFFFF187FF;
defparam sdpb_inst_5.INIT_RAM_39 = 256'hA01BDDEFFFFFFFFF02FF04FFFFF83CBFFFFFF861202800BF9DFFFFFFFFE08FF8;
defparam sdpb_inst_5.INIT_RAM_3A = 256'hFFFFF1193FFFFFFE0C0F08817F8F7FFFFFFFF841C19FFFFF0383FFFFFFC386C0;
defparam sdpb_inst_5.INIT_RAM_3B = 256'h34FF1FDFFFFFFFFF8060FFFFFF5003FFFFFFF03014BC27F8FBFFFFFFFFF0E263;
defparam sdpb_inst_5.INIT_RAM_3C = 256'hFFFCA053FFFFFFFC0689029FF1FFFFFFFFFFFF007FFFFFC2053FFFFFFF819070;
defparam sdpb_inst_5.INIT_RAM_3D = 256'h4FE3FCFFFFFFFFFFFFFFFFFFE0003FFFFFFFF0186809FE1FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3E = 256'hFFFFC47FFFFFFFFF008EC27E3FFFFFFFFFFFFFFFFFFFFF1C27FFFFFFFFC021B0;
defparam sdpb_inst_5.INIT_RAM_3F = 256'hBCFFEFFFFFFFFFFFFFFFFFFFFF1FFFFFFFFFFE023B13E7FFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[6]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b1;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'h8002D3AF8830000000000000000000002FFFFFFF00000048C302400000000002;
defparam sdpb_inst_6.INIT_RAM_01 = 256'h0000000001FFFFBFFFF28405EFFEFEE60800000000000000000002FF6FFFF580;
defparam sdpb_inst_6.INIT_RAM_02 = 256'hF7FFFFFBB7000000000000000000003FFBFDFFEDB1B8FFFFFCF9F80000000000;
defparam sdpb_inst_6.INIT_RAM_03 = 256'h00000000FFBC67EBEE80AFFFFFFFD7320000000000000000002BFE1F9BFFFC05;
defparam sdpb_inst_6.INIT_RAM_04 = 256'hFFF4DFFE7086000000000000000003F7F8FF0028125FF7FFFFFB040000000000;
defparam sdpb_inst_6.INIT_RAM_05 = 256'h00000007E3C799FC00007FFFFFFFF8040000000000000000005EFF07E700012F;
defparam sdpb_inst_6.INIT_RAM_06 = 256'h9D9FF9FD102002000000000000048F81FE3FE0000FF83FFE7FE1C80000000000;
defparam sdpb_inst_6.INIT_RAM_07 = 256'h0000033FC8F9E300002FE68CEFFFF002000000000000000003FE3FC0F80002FF;
defparam sdpb_inst_6.INIT_RAM_08 = 256'hC01FFFFC5004A000000000000004F1E23F800002FCE383FFFF84020000000000;
defparam sdpb_inst_6.INIT_RAM_09 = 256'h0000044FF03F000009FC2000FFFFB9000000000000000000007F8FF800009B47;
defparam sdpb_inst_6.INIT_RAM_0A = 256'h6F1FDDD1400192000000000000203E78C0200037C105C7FB7BE1080120000000;
defparam sdpb_inst_6.INIT_RAM_0B = 256'h00001003FE00000000407F79FFFFA0100161000000000000348FE00200009601;
defparam sdpb_inst_6.INIT_RAM_0C = 256'h9E7FFFC4808240000000000000008FC62000000001FBCFFFF7AA73C408000000;
defparam sdpb_inst_6.INIT_RAM_0D = 256'h000082040501000000005DF1FFF5E2029480000000000000013A02000000840F;
defparam sdpb_inst_6.INIT_RAM_0E = 256'h7C3FFA880746400000000000004A0800400000E003EF8FFFF0412AA000000000;
defparam sdpb_inst_6.INIT_RAM_0F = 256'h010400910080000000807BC09FD003BF0000000000000048200000000440400F;
defparam sdpb_inst_6.INIT_RAM_10 = 256'hF01540001F90000000401000000010580009000403DE81F45110BD4000000080;
defparam sdpb_inst_6.INIT_RAM_11 = 256'h80000002000000000100FC000020A4970000000020000043002180000000201E;
defparam sdpb_inst_6.INIT_RAM_12 = 256'h0000008E16000000000000006004100000000000070000410104C50000000031;
defparam sdpb_inst_6.INIT_RAM_13 = 256'h00042A0000000000000200000009614E00000008000000100000000800000030;
defparam sdpb_inst_6.INIT_RAM_14 = 256'h00000261F8000000000010001081000004000040000000001ABA900000000002;
defparam sdpb_inst_6.INIT_RAM_15 = 256'h0000400000020000002000020048726000000008000000462000002000000100;
defparam sdpb_inst_6.INIT_RAM_16 = 256'h00000191000000000000000000000000100020010000000063A8000000000008;
defparam sdpb_inst_6.INIT_RAM_17 = 256'h0000000000020C0000C000000010380000000080080000000000008098001800;
defparam sdpb_inst_6.INIT_RAM_18 = 256'hE00083F100000000403C00000000000000800006000000062DC0000000000080;
defparam sdpb_inst_6.INIT_RAM_19 = 256'h000000000000002000F0FD0000EB8000000000FE800000000000000001001001;
defparam sdpb_inst_6.INIT_RAM_1A = 256'hC1022F80000000002F00000000000000000040006F780833220000000001B800;
defparam sdpb_inst_6.INIT_RAM_1B = 256'h0000000000000000001F7C0417700000000000000000000000000000120003BD;
defparam sdpb_inst_6.INIT_RAM_1C = 256'h081B18000000000000000000000000001A000000F8E000C50000000000000000;
defparam sdpb_inst_6.INIT_RAM_1D = 256'h00800007E0000000003B9800152000000000000A8000000000007800000007E6;
defparam sdpb_inst_6.INIT_RAM_1E = 256'h0096C00000000000148000000006000000000001CEC000300000000000037800;
defparam sdpb_inst_6.INIT_RAM_1F = 256'h0003000021000300007E60026200000000000690000010070000000020800F9E;
defparam sdpb_inst_6.INIT_RAM_20 = 256'h10C000000000000040000020C000100000000003FB8000400000000000100000;
defparam sdpb_inst_6.INIT_RAM_21 = 256'h880010000000000200F5E0014000000000010800000420001000000000081CEC;
defparam sdpb_inst_6.INIT_RAM_22 = 256'h1000000000000020000023000200000000000007E60000000000000001000000;
defparam sdpb_inst_6.INIT_RAM_23 = 256'h008000000000000001EEE0020000000000020000084000800000000005003F98;
defparam sdpb_inst_6.INIT_RAM_24 = 256'h00000000000108000001000000000000000000075F0000000000000040000008;
defparam sdpb_inst_6.INIT_RAM_25 = 256'h00000000000000000199C0000000000001800000200000000000000000003E68;
defparam sdpb_inst_6.INIT_RAM_26 = 256'h00000000000A000000400000000000000000000E360000000000001000000000;
defparam sdpb_inst_6.INIT_RAM_27 = 256'h000000000000000003F780000000000840000008000000000000000000007ED0;
defparam sdpb_inst_6.INIT_RAM_28 = 256'h0000000022800000200000000000000000000019EC00000000000C0000010020;
defparam sdpb_inst_6.INIT_RAM_29 = 256'h000000000000000003EF00000000E51000000200000000000000000000007560;
defparam sdpb_inst_6.INIT_RAM_2A = 256'h00000FE0A0000004010000000000000000000013D80000007F03000000400000;
defparam sdpb_inst_6.INIT_RAM_2B = 256'h000000000000000007DC000001FE4F000000800000000000000000000000EAC0;
defparam sdpb_inst_6.INIT_RAM_2C = 256'h0003E03FC000010000000000000000000000002BB800003F01F8000008000000;
defparam sdpb_inst_6.INIT_RAM_2D = 256'h0003F000000000000FBC00003C01F8000010000000000018000000000003D580;
defparam sdpb_inst_6.INIT_RAM_2E = 256'h00EC0BF400002008000000027FC0000000000057C00005C01F80000200000000;
defparam sdpb_inst_6.INIT_RAM_2F = 256'h0BFFFC00000000001FC0002FE07E40000200000000007FFF000000000003FC00;
defparam sdpb_inst_6.INIT_RAM_30 = 256'h3FFFF900000400000000017FF7E00000000000F80008BF9FC800000010000000;
defparam sdpb_inst_6.INIT_RAM_31 = 256'hFE07C6000000000000007C7FFF60000040000000002FF1DD8000000000000003;
defparam sdpb_inst_6.INIT_RAM_32 = 256'h3F2EC0000040100000005FC01E180000000000000F87EFEC0000040000000003;
defparam sdpb_inst_6.INIT_RAM_33 = 256'h8001E50000000000000CC160E80000080000000009F8007800000000000001F0;
defparam sdpb_inst_6.INIT_RAM_34 = 256'h00E80000080000000013F0003FAC0000000000001BC00E80000000000000009E;
defparam sdpb_inst_6.INIT_RAM_35 = 256'h007FFA900000000004001E0680000080200000003BC007FFB0000000000001FF;
defparam sdpb_inst_6.INIT_RAM_36 = 256'h018000010000000001F792010FF0000000000000000028000008000000001F36;
defparam sdpb_inst_6.INIT_RAM_37 = 256'h2200C0F00000000000000110000010040000001FFF49000C6000000000000000;
defparam sdpb_inst_6.INIT_RAM_38 = 256'h20000010000000000F7FEEC00C0380000000000000230000010000000001FFFF;
defparam sdpb_inst_6.INIT_RAM_39 = 256'hA01821F00000000011340C00000000800000006BF02800801E0000000004700C;
defparam sdpb_inst_6.INIT_RAM_3A = 256'h00000101000000000F7E0081001F800000000060018000001000000000032F80;
defparam sdpb_inst_6.INIT_RAM_3B = 256'h34000FC00000000000600000001010000000003FF8042001FC00000000009CE0;
defparam sdpb_inst_6.INIT_RAM_3C = 256'h0000A01000000000077F018001FE00000000000000000000050000000001FFC0;
defparam sdpb_inst_6.INIT_RAM_3D = 256'h4003FF000000000000000000000000000000001FFA00001F7000000000000000;
defparam sdpb_inst_6.INIT_RAM_3E = 256'h000004000000000000FFC2003FF0000000000000000000000000000000003FF0;
defparam sdpb_inst_6.INIT_RAM_3F = 256'h80FFE00000000000000000000000000000000003FF1007FF0000000000000000;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[7]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b1;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFF;
defparam sdpb_inst_7.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC03FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_03 = 256'hFFFFFFFFFFC3981FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE067FFFFFF;
defparam sdpb_inst_7.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80700FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_05 = 256'hFFFFFFFF9C386603FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00F818FFFFFF;
defparam sdpb_inst_7.INIT_RAM_06 = 256'hE07FFFFFFFFFFFFFFFFFFFFFFFFFF07E01C01FFFFFFFCFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_07 = 256'hFFFFFFC037061CCFFFFFF873FFFFFFFFFFFFFFFFFFFFFFFFFC01C03F06FFFFFF;
defparam sdpb_inst_7.INIT_RAM_08 = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFB0E1DC070FFFFFF1C0FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_09 = 256'hFFFFFC300FC0D0FFFFFFC007FFFFFFFFFFFFFFFFFFFFFFFFCF8070070FFFFFF8;
defparam sdpb_inst_7.INIT_RAM_0A = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFC3C187311FFFFFFE003FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0B = 256'hFFFFE91C01C18FFFFFFF8007FFFFFFFFFFFFFFFFFFFFFFFE03701E14FFFFFFF0;
defparam sdpb_inst_7.INIT_RAM_0C = 256'h01FFFFFFFFFFFFFFFFFFFFFFFF70703010FFFFFFFE003FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0D = 256'hFFFF0C438290FFFE000F800FFFFFFFFFFFFFFFFFFFFFFFF184C4650FFFFC13F0;
defparam sdpb_inst_7.INIT_RAM_0E = 256'h03FFFFFFFFFFFFFFFFFFFFFFF89410310FFFC0001C007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0F = 256'h38F9C308A10FFF8FFF07801FFFFFFFFFFFFFFFFFFFE3FFA4418618FFF83F81F0;
defparam sdpb_inst_7.INIT_RAM_10 = 256'h000FFFFFFFFFFFFFFFB0E38FC62CA201FFF0FFF83C007FFFFFFFFFFFFFFFFF0E;
defparam sdpb_inst_7.INIT_RAM_11 = 256'h3FF270810FFFF1FFFE1F00003FFFFFFFFFFFFFF1C739FC383C083FFF1FFFC3E0;
defparam sdpb_inst_7.INIT_RAM_12 = 256'h0007FFFFFFFFFFFFFE0003FF810861FFFF1FFFF1F80000FFFFFFFFFFFFFF0600;
defparam sdpb_inst_7.INIT_RAM_13 = 256'hFFF89517FFFF8FFFE1FC00003FFFFFFFFFFFFFF0003FFF0CC93FFFF0FFFF1FC0;
defparam sdpb_inst_7.INIT_RAM_14 = 256'h003FFFFFFFFFFFFFFF800FFFE860FFFFF87FFC3FE00003FFFFFFFFFFFFFFC001;
defparam sdpb_inst_7.INIT_RAM_15 = 256'hFFFE27FFFFFC1FE0FFC00001FFFFFFFFFFFFFFF000FFFF801FFFFFC3FF87FE00;
defparam sdpb_inst_7.INIT_RAM_16 = 256'h03FFFFFFFFFFFFFFF0007FFFFAFFFFFFE0401FFE00003FFFFFFFFFFFFFFF0007;
defparam sdpb_inst_7.INIT_RAM_17 = 256'hFFFFFFFFFFFC03FFFF00003FFFFFFFFFFFFFFF0007FFFFFFFFFFFF0007FFE000;
defparam sdpb_inst_7.INIT_RAM_18 = 256'h1FFFFFFFFFFFFFFF8003FFFFFFFFFFFFFF7FFFF80003FFFFFFFFFFFFFFF8007F;
defparam sdpb_inst_7.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFF007FFFFFFFFFFFFFFFFFFFE000;
defparam sdpb_inst_7.INIT_RAM_1A = 256'h3FFFFFFFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFFFF8007FFFFFFFFFFFFFFFE07FF;
defparam sdpb_inst_7.INIT_RAM_1B = 256'hFFFFFFFFFFFF83FFFFE003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_7.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFF3FFFFFFFFFFFFFE1FFFFFF001FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1D = 256'hC07FFFF81FFFFFFFFFC007FFFFFFFFFFFFFFFFE07FFFFFFFFFFF87FFFFFFF800;
defparam sdpb_inst_7.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFC07FF801FFF9FFFFFFFFFFFE003FFFFFFFFFFFFFFFFC07FF;
defparam sdpb_inst_7.INIT_RAM_1F = 256'h01FCFFFFC00000FFFF800FFFFFFFFFFFFFFFF80FFF800FF8FFFFFFFFCFFFF001;
defparam sdpb_inst_7.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFF03FFF801F3FFF8FFFFFFFFFFC007FFFFFFFFFFFFFFF81FFF8;
defparam sdpb_inst_7.INIT_RAM_21 = 256'h77FFE7FFFFFFFFFFFF001FFFFFFFFFFFFFFE07FFFC03DFFFCFFFFFFFFFFFE003;
defparam sdpb_inst_7.INIT_RAM_22 = 256'hFFFFFFFFFFFFFC1FFFFE1CFFF9FFFFFFFFFFFFF800FFFFFFFFFFFFFFE0FFFFC0;
defparam sdpb_inst_7.INIT_RAM_23 = 256'hFF3FFFFFFFFFFFFFFE001FFFFFFFFFFFFF81FFFFF7BFFE7FFFFFFFFFFFFFC007;
defparam sdpb_inst_7.INIT_RAM_24 = 256'hFFFFFFFFFFFE07FFFFFEFFEFFFFFFFFFFFFFFFF800FFFFFFFFFFFFF03FFFFFF7;
defparam sdpb_inst_7.INIT_RAM_25 = 256'h7FFFFFFFFFFFFFFFFE003FFFFFFFFFFFE07FFFFFDFFBFFFFFFFFFFFFFFFFC007;
defparam sdpb_inst_7.INIT_RAM_26 = 256'hFFFFFFFFFF81FFFFFFBFEFFFFFFFFFFFFFFFFFF001FFFFFFFFFFFC0FFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFC007FFFFFFFFFF03FFFFFF7FDFFFFFFFFFFFFFFFFFF800F;
defparam sdpb_inst_7.INIT_RAM_28 = 256'hFFFFFFFFC07FFFFFDFFBFFFFFFFFFFFFFFFFFFE003FFFFFFFFFE03FFFFFEFFDF;
defparam sdpb_inst_7.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFF800FFFFFFFF180FFFFFFDFF7FFFFFFFFFFFFFFFFFFF001F;
defparam sdpb_inst_7.INIT_RAM_2A = 256'hFFFFF0001FFFFFFBFEFFFFFFFFFFFFFFFFFFFFC007FFFFFF8000FFFFFFBFEFFF;
defparam sdpb_inst_7.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFF001FFFFFE0000FFFFFF7FDFFFFFFFFFFFFFFFFFFFFE003F;
defparam sdpb_inst_7.INIT_RAM_2C = 256'hFFFC00003FFFFEFFBFFFFFFFFFFFFFFFFFFFFF8007FFFFC00007FFFFF7FFFFFF;
defparam sdpb_inst_7.INIT_RAM_2D = 256'hFFF00FFFFFFFFFFFE003FFFFC00003FFFFEFFFFFFFFFFFC7FFFFFFFFFFFC007F;
defparam sdpb_inst_7.INIT_RAM_2E = 256'hFF000003FFFFDFF7FFFFFFFC003FFFFFFFFFFF003FFFF800003FFFFDFF7FFFFF;
defparam sdpb_inst_7.INIT_RAM_2F = 256'hF00003FFFFFFFFFFC03FFFD000003FFFFDFFFFFFFFFF8000FFFFFFFFFFF803FF;
defparam sdpb_inst_7.INIT_RAM_30 = 256'hC00000FFFFFBFEFFFFFFFE00081FFFFFFFFFFF07FFF7400007FFFFFFEFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_31 = 256'h000001FFFFFFFFFFFFFF8000001FFFFFBFEFFFFFFFC000207FFFFFFFFFFFFFFC;
defparam sdpb_inst_7.INIT_RAM_32 = 256'h00003FFFFFBFEFFFFFFF80000007FFFFFFFFFFFFF0000003FFFFFBFEFFFFFFFC;
defparam sdpb_inst_7.INIT_RAM_33 = 256'h000000FFFFFFFFFFFFC0000007FFFFF7FFFFFFFFF00000003FFFFFFFFFFFFE00;
defparam sdpb_inst_7.INIT_RAM_34 = 256'h0007FFFFF7FDFFFFFFE000000003FFFFFFFFFFFC0000007FFFFF7FDFFFFFFF01;
defparam sdpb_inst_7.INIT_RAM_35 = 256'h0000006FFFFFFFFFF80000007FFFFF7FDFFFFFFE040000000FFFFFFFFFFFC000;
defparam sdpb_inst_7.INIT_RAM_36 = 256'h007FFFFEFFBFFFFFFE086C0EF000FFFFFFFFFFC0000007FFFFF7FBFFFFFFE0C9;
defparam sdpb_inst_7.INIT_RAM_37 = 256'hDDFF000FFFFFFFFFE000000FFFFFEFFBFFFFFFE000B0FFF007FFFFFFFFFC0000;
defparam sdpb_inst_7.INIT_RAM_38 = 256'h1FFFFFEFF7FFFFFFF000013FF0007FFFFFFFFF000000FFFFFEFF7FFFFFFE0000;
defparam sdpb_inst_7.INIT_RAM_39 = 256'h5FE0000FFFFFFFFFE00003FFFFFCFF7FFFFFFF800017FF0001FFFFFFFFF80000;
defparam sdpb_inst_7.INIT_RAM_3A = 256'hFFFFF8FEFFFFFFFFF000017E00007FFFFFFFFF80007FFFFFCFEFFFFFFFFC0000;
defparam sdpb_inst_7.INIT_RAM_3B = 256'h0800003FFFFFFFFFFF9FFFFFFF8FCFFFFFFFFFC00003C00003FFFFFFFFFF001F;
defparam sdpb_inst_7.INIT_RAM_3C = 256'hFFFF1F8FFFFFFFFFF80000000001FFFFFFFFFFFFFFFFFFF9F8FFFFFFFFFE0000;
defparam sdpb_inst_7.INIT_RAM_3D = 256'h000000FFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFE0040000000FFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3E = 256'hFFFFFBFFFFFFFFFFFF000000000FFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFFC000;
defparam sdpb_inst_7.INIT_RAM_3F = 256'h00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000FFFFFFFFFFFFFFFF;

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[23:0],sdpb_inst_8_dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_1}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_8.READ_MODE = 1'b1;
defparam sdpb_inst_8.BIT_WIDTH_0 = 8;
defparam sdpb_inst_8.BIT_WIDTH_1 = 8;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_8.RESET_MODE = "SYNC";
defparam sdpb_inst_8.INIT_RAM_00 = 256'hA3A2A3A3A4A3A3A3A3A2A2A2A2A0A09D9A9691887357534F6465625B61450B15;
defparam sdpb_inst_8.INIT_RAM_01 = 256'hA1A2A2A2A3A2A3A2A2A2A2A3A1A3A2A2A2A2A1A2A2A2A3A4A2A3A3A4A4A4A4A3;
defparam sdpb_inst_8.INIT_RAM_02 = 256'hA2A3A2A3A1A3A2A1A3A1A0A2A2A2A2A3A1A2A1A0A1A0A1A1A0A1A0A1A1A0A1A0;
defparam sdpb_inst_8.INIT_RAM_03 = 256'hA7A6A7A6A4A4A5A5A4A5A6A7A5A5A5A5A5A5A4A5A5A5A6A4A3A4A4A4A2A4A4A2;
defparam sdpb_inst_8.INIT_RAM_04 = 256'h747571736C6B62A1A2A4A6A7A7A8A8A9A7A8A7A7A8A7A8A8A7A7A7A7A6A6A4A5;
defparam sdpb_inst_8.INIT_RAM_05 = 256'hA3A1A2A09F9D9B9790836F53545D64625E2E181010520E1412140C7567757574;
defparam sdpb_inst_8.INIT_RAM_06 = 256'hA1A0A1A2A2A1A2A1A1A1A2A1A2A1A2A2A1A3A2A2A2A3A3A3A3A4A4A5A4A3A3A3;
defparam sdpb_inst_8.INIT_RAM_07 = 256'hA1A1A1A1A0A0A1A1A1A0A19FA0A0A1A0A1A1A1A1A0A1A2A2A1A1A2A0A1A1A3A0;
defparam sdpb_inst_8.INIT_RAM_08 = 256'hA5A5A4A3A4A4A4A4A5A5A6A4A3A4A4A3A4A2A2A2A1A2A2A1A1A0A1A0A1A0A1A1;
defparam sdpb_inst_8.INIT_RAM_09 = 256'hA6A7A7A7A6A7A6A6A7A7A6A8A6A5A6A5A5A6A5A6A5A6A4A5A5A5A3A4A4A5A4A5;
defparam sdpb_inst_8.INIT_RAM_0A = 256'h6A525364654C3B54643C10175D7372737562757574747370626F7D9FA2A5A6A6;
defparam sdpb_inst_8.INIT_RAM_0B = 256'hA1A1A0A1A2A3A2A2A1A2A1A2A2A2A4A4A4A5A4A4A4A4A4A3A2A19F9C99948F81;
defparam sdpb_inst_8.INIT_RAM_0C = 256'h9F9F9F9FA0A0A1A0A1A1A09FA2A1A1A0A0A0A1A0A1A1A1A0A0A1A0A09FA0A1A1;
defparam sdpb_inst_8.INIT_RAM_0D = 256'hA4A3A4A3A4A2A2A1A19FA0A0A09F9F9E9EA0A0A0A19FA0A0A0A09FA0A1A0A0A1;
defparam sdpb_inst_8.INIT_RAM_0E = 256'hA7A4A6A5A5A4A3A5A5A4A5A4A4A4A3A3A4A2A3A3A5A4A4A4A5A3A3A5A4A4A4A3;
defparam sdpb_inst_8.INIT_RAM_0F = 256'h7A76757674735F7373736F706D599CA1A1A4A5A7A6A6A5A7A5A5A6A6A5A5A7A4;
defparam sdpb_inst_8.INIT_RAM_10 = 256'hA3A2A4A5A4A5A4A6A4A6A6A4A4A2A3A09F9A97938A7F69574E625D6255636D82;
defparam sdpb_inst_8.INIT_RAM_11 = 256'h9F9FA19F9F9FA09E9F9EA09FA0A09EA0A09F9FA0A19E9FA0A1A1A2A1A3A1A1A2;
defparam sdpb_inst_8.INIT_RAM_12 = 256'h9FA09F9F9E9F9EA09EA09E9FA09FA09EA09F9D9F9FA09F9F9F9EA0A0A09E9FA0;
defparam sdpb_inst_8.INIT_RAM_13 = 256'hA3A3A1A3A5A2A3A2A3A4A4A3A3A2A3A1A3A2A3A2A4A3A3A2A4A1A09FA09EA0A0;
defparam sdpb_inst_8.INIT_RAM_14 = 256'h757C9DA2A4A3A4A5A6A6A6A6A7A6A4A5A5A5A5A7A5A5A3A3A2A3A3A3A5A2A3A2;
defparam sdpb_inst_8.INIT_RAM_15 = 256'hA4A5A3A4A2A09E9A959287786B5858052A5855617A757576777374547272706F;
defparam sdpb_inst_8.INIT_RAM_16 = 256'h9E9E9E9E9E9E9E9F9E9E9F9E9F9F9EA09FA0A1A1A1A2A2A3A4A4A4A5A4A5A6A4;
defparam sdpb_inst_8.INIT_RAM_17 = 256'h9D9D9EA09E9E9E9E9F9E9F9F9F9E9F9E9F9F9E9E9E9F9D9E9E9F9E9F9D9E9E9E;
defparam sdpb_inst_8.INIT_RAM_18 = 256'hA2A2A2A0A3A3A2A2A2A1A2A2A1A09F9F9F9C9D9F9F9E9D9E9D9D9D9E9D9C9D9E;
defparam sdpb_inst_8.INIT_RAM_19 = 256'hA4A5A3A5A5A6A6A4A3A3A2A1A1A2A0A2A2A2A2A2A1A1A1A1A0A0A2A2A0A2A1A2;
defparam sdpb_inst_8.INIT_RAM_1A = 256'h83796E4E0B694B595A6472757165308463716D65569A9EA1A3A5A4A5A4A4A5A2;
defparam sdpb_inst_8.INIT_RAM_1B = 256'h9F9E9D9E9FA1A1A1A1A1A1A3A3A4A3A5A4A5A7A6A7A6A5A5A4A3A39F9D9A948E;
defparam sdpb_inst_8.INIT_RAM_1C = 256'h9D9E9D9D9E9E9D9D9E9C9B9D9E9D9D9D9E9D9D9D9D9D9C9F9D9D9D9D9D9D9E9C;
defparam sdpb_inst_8.INIT_RAM_1D = 256'hA09E9E9D9C9D9E9E9D9D9D9B9E9C9D9C9E9C9B9C9D9E9C9D9D9C9D9D9B9D9D9D;
defparam sdpb_inst_8.INIT_RAM_1E = 256'hA2A0A0A1A0A1A1A1A29FA0A19FA2A0A19FA0A1A0A0A1A1A09FA1A0A2A2A09FA1;
defparam sdpb_inst_8.INIT_RAM_1F = 256'h0C7D7C787569625F959EA0A2A3A4A3A4A4A4A5A4A5A5A2A4A5A5A3A4A3A3A2A2;
defparam sdpb_inst_8.INIT_RAM_20 = 256'hA3A3A3A4A5A5A6A6A6A6A6A6A5A4A4A2A29F9C98938C867D704D1055295F8B69;
defparam sdpb_inst_8.INIT_RAM_21 = 256'h9B9D9C9B9D9B9C9C9C9B9A9B9B9B9C9C9C9D9C9C9D9D9E9D9E9F9FA1A0A0A1A2;
defparam sdpb_inst_8.INIT_RAM_22 = 256'h9B9C9B9B9A9B9B9C9B9C9B9A9C9D9D9E9C9C9C9D9C9D9C9C9C9C9C9C9C9C9C9D;
defparam sdpb_inst_8.INIT_RAM_23 = 256'hA0A0A09F9F9FA09FA0A09F9F9EA09FA1A0A0A09D9E9D9E9D9C9C9C9D9B9B9A9B;
defparam sdpb_inst_8.INIT_RAM_24 = 256'hA4A4A5A4A4A4A2A3A4A6A2A4A3A3A4A3A2A2A2A1A0A09E9E9F9EA0A0A19F9F9E;
defparam sdpb_inst_8.INIT_RAM_25 = 256'hA7A6A6A5A3A3A09E9C98938E877B6A544F4361847F7A0F70776961939B9FA1A2;
defparam sdpb_inst_8.INIT_RAM_26 = 256'h9B9A9B9B9B9A9C9B9C9C9B9E9E9E9DA09E9FA0A1A1A3A2A2A4A4A5A5A6A6A6A6;
defparam sdpb_inst_8.INIT_RAM_27 = 256'h9A9B9B9B9B9B9B9C9B9B9A9C9B9B9D9B9C9C9B9B9C9C9A9A9A9A9A9C9A999B9A;
defparam sdpb_inst_8.INIT_RAM_28 = 256'h9D9E9E9F9F9E9F9E9D9C9C9B9B9C9C9B9C99999C9A9A9A999B9A9A999B9A999A;
defparam sdpb_inst_8.INIT_RAM_29 = 256'hA2A2A3A19FA1A1A1A0A09D9D9F9D9F9E9E9F9E9E9E9F9F9E9F9FA09F9E9D9F9F;
defparam sdpb_inst_8.INIT_RAM_2A = 256'h9691897D736A6A72716E7385545697989DA1A1A3A3A3A3A4A2A5A2A2A2A1A3A3;
defparam sdpb_inst_8.INIT_RAM_2B = 256'h9D9C9E9E9E9FA0A0A1A2A2A2A1A2A4A4A5A4A7A6A5A6A7A6A5A4A3A29F9F9D98;
defparam sdpb_inst_8.INIT_RAM_2C = 256'h9B99999B9A9A999A9A9B9A9A99999B9A999A9A9A999A9A9B9B989B9A9B9C9B9B;
defparam sdpb_inst_8.INIT_RAM_2D = 256'h99989A9A9A9A9B9999989799989A9A9A9A9A9999999A9A99999A9999999B9A9C;
defparam sdpb_inst_8.INIT_RAM_2E = 256'h9C9C9D9D9E9E9C9F9E9D9E9C9C9C9C9C9D9C9D9E9B9E9E9C9C9C9B999B9B9C9B;
defparam sdpb_inst_8.INIT_RAM_2F = 256'h91969C9EA0A1A2A3A3A4A2A4A3A3A3A3A2A1A2A3A09FA1A1A2A0A09F9D9E9D9C;
defparam sdpb_inst_8.INIT_RAM_30 = 256'hA2A1A3A4A5A5A6A5A6A6A6A6A6A5A5A4A5A3A2A19F9B9895938F898383858A8D;
defparam sdpb_inst_8.INIT_RAM_31 = 256'h9899989898999796989798989A989898969899999A9B9B9D9C9D9D9E9F9FA0A1;
defparam sdpb_inst_8.INIT_RAM_32 = 256'h969598969898979B989998999799989A9998979899989899999A989898989898;
defparam sdpb_inst_8.INIT_RAM_33 = 256'h9C9C9C9C9B9B9C9D9B9A9B9B9B9A9A9A9B989898979997979896979898989996;
defparam sdpb_inst_8.INIT_RAM_34 = 256'hA3A3A3A2A1A2A0A1A0A3A1A19E9F9E9F9D9C9D9C9C9B9C9B9D9D9C9C9E9D9C9C;
defparam sdpb_inst_8.INIT_RAM_35 = 256'hA5A5A6A5A5A4A4A3A0A29F9D9C9B9A999994989B9A9D9FA0A1A3A4A3A2A4A2A3;
defparam sdpb_inst_8.INIT_RAM_36 = 256'h9596969697979897989A9999999C9D9C9DA09EA0A1A0A3A2A2A4A4A5A5A4A5A6;
defparam sdpb_inst_8.INIT_RAM_37 = 256'h9897979798969698969697979999989997969798979597969797959796979597;
defparam sdpb_inst_8.INIT_RAM_38 = 256'h9997989698969797949698979596949696979797969596989697979595979698;
defparam sdpb_inst_8.INIT_RAM_39 = 256'h000000000000009A98999A9A9A9B9C9B9B9A9A9B9B9B9A989C999A9A999A9998;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clkb),
  .CE(oce)
);
MUX2 mux_inst_6 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_8_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(dout[1]),
  .I0(sdpb_inst_1_dout[1]),
  .I1(sdpb_inst_8_dout[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_20 (
  .O(dout[2]),
  .I0(sdpb_inst_2_dout[2]),
  .I1(sdpb_inst_8_dout[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_27 (
  .O(dout[3]),
  .I0(sdpb_inst_3_dout[3]),
  .I1(sdpb_inst_8_dout[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_34 (
  .O(dout[4]),
  .I0(sdpb_inst_4_dout[4]),
  .I1(sdpb_inst_8_dout[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_41 (
  .O(dout[5]),
  .I0(sdpb_inst_5_dout[5]),
  .I1(sdpb_inst_8_dout[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_48 (
  .O(dout[6]),
  .I0(sdpb_inst_6_dout[6]),
  .I1(sdpb_inst_8_dout[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_55 (
  .O(dout[7]),
  .I0(sdpb_inst_7_dout[7]),
  .I1(sdpb_inst_8_dout[7]),
  .S0(dff_q_1)
);
endmodule //Gowin_SDPB4
