//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Tue Sep 05 13:32:03 2023

module Gowin_SDPB3 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);//gaussian_blur_3x3 - new

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [15:0] ada;
input [7:0] din;
input [15:0] adb;

wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [0:0] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [1:1] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [1:1] sdpb_inst_3_dout;
wire [29:0] sdpb_inst_4_dout_w;
wire [1:0] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [2:2] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [2:2] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [3:3] sdpb_inst_7_dout;
wire [30:0] sdpb_inst_8_dout_w;
wire [3:3] sdpb_inst_8_dout;
wire [29:0] sdpb_inst_9_dout_w;
wire [3:2] sdpb_inst_9_dout;
wire [30:0] sdpb_inst_10_dout_w;
wire [4:4] sdpb_inst_10_dout;
wire [30:0] sdpb_inst_11_dout_w;
wire [4:4] sdpb_inst_11_dout;
wire [30:0] sdpb_inst_12_dout_w;
wire [5:5] sdpb_inst_12_dout;
wire [30:0] sdpb_inst_13_dout_w;
wire [5:5] sdpb_inst_13_dout;
wire [29:0] sdpb_inst_14_dout_w;
wire [5:4] sdpb_inst_14_dout;
wire [30:0] sdpb_inst_15_dout_w;
wire [6:6] sdpb_inst_15_dout;
wire [30:0] sdpb_inst_16_dout_w;
wire [6:6] sdpb_inst_16_dout;
wire [30:0] sdpb_inst_17_dout_w;
wire [7:7] sdpb_inst_17_dout;
wire [30:0] sdpb_inst_18_dout_w;
wire [7:7] sdpb_inst_18_dout;
wire [29:0] sdpb_inst_19_dout_w;
wire [7:6] sdpb_inst_19_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_3;
wire mux_o_9;
wire mux_o_15;
wire mux_o_21;
wire mux_o_27;
wire mux_o_33;
wire mux_o_39;
wire mux_o_45;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b1;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h1832D9F2094634DC0722DBFEA77A12E4A85C80FCDE1FDDE9F7F3A238FBCA1DFC;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hDF97C54923E7976EBFAE764982136BAFCC39B6CFBEFB6FE38710EE8A0E73AD25;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h542C8950A92E0393F27D8FBA46002E029F7DBCAF7B860C03C5CF71F57AC73362;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h39754F84E0F484298F121DE61E500404E37CB7EA828E8804861CF19D6555855C;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h2F02F01C687E41501EBF85EF86D40003D002F0DC904651AE11C4407A118FBECD;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hE92824F2F0E985562DB42E10E185DF00BD20772B00B815FC6135401F401021EB;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hF0E5DC1D48E1194FF9D82F1125A0F92E4790473A1865075D5FA03806E4348E16;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h7FDCF21686418DD22FCBA7F8308560D19D240DB79A0F1073FBF5906E4A5A80F7;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h0B536B80CA8F7BB2D3F8C67E83C0D8C325815C16BE50F0040A17B4243369C650;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h59ED831E8D8D761B921C3DB77420038767187AE9FB7B060C61E9BA0C008CFAE1;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h9BB80ACFDFA2F6A9501CAFF0BE450E06F901CEEDB47EB5F0740B56CEC93375F9;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h3FF3C6266B22987480C86CDFE5A807651CDAB015E588E58300000377D0AFA903;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h51066F011DBAAEE0E84437D6BCBF267DFE6C585DECBC8050000000B78EC66EA0;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hC7DD80D810DA0394C11DE3E9A3EB5C69F242A1607104B0FE00000411A9E1207D;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h49CF696CBC93B85F2DA8C37C3ED0A34A5C3F1DA806750BBFE37034CD7AEA544F;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hA5CBD7334E294675BE4D33DBF85581AD0F1C7065FB889F47FA4F056C5883B023;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h20CE067296DB282B779532A4F0DC5F04D7FB43582FDA1CBE07031140C307F101;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h08077FFB9ADBC5F8256DA5DD8B87A39FE979B1FB484C1AC7FDB45E116F0B3DAC;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h57600AFFF3CDEFFC08FDD733A77CC60EA02C734F0B90BBE3AFE13378F8D730BF;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h8371481B95DEBBD6942B705A784B93EF98A5A24AA4F74C548F0570FEC160A58A;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h23638E817E7F5FF77B96F7A48213E826DF0FED3F7C21D01F23CC2595ACA34684;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hA6C29F14001E657EDCF20D798237871432F20D1594441683FE02391202C8EF8F;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h376A9B040C17BFFE1C8F532AFA146382C327B0245853561A128489A380065B03;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h30A39D7DE8C7BFFBF3787FCC4D07DF7E45A1F0FDD87CC235E3945842FE515675;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h10A53AFBFEC406F9C7A38DF72EFDB4F063013737C08D65B4A618C95827750E02;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h47A50D5B5D45BC536F66E145767C6F37D9407FFF7E90C0D861FA13E6103EFEFF;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hBEB0A25B56BFF943F75DC374ECB8A2367A8A11F9FF208B046B1DBAFD0BDDD30B;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h4E71A0B6EC7F9EC0FBFCEC32A26E340E50C808278CCE4318192410919BA8DD85;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h59FC2C42C2A1DECB8FF5FFE736F539980CDF0BE5BF75B1277382BD4D96B2658F;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hD2A8CC70B86B8CFEE0FFBB3F19FB0B323337122E63FFDD5EB7DA1344134453BE;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h385A5782D4C65437FE239BFFC37CF1814775BFBABE8720925EC5EA62C0E13765;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hEF4608487A5119566F8279B3F80B14C5DCBF371D7FF320040C27C88342F26C32;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h150231806C710428A0D0AC97A3C4E2FD8B935B7F90B6DA16539C5FDF07075B5A;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h211430A84B6EBD611C6881EFF4ED2F34F5448AB1E72CB0B4BCB904952378B0BF;
defparam sdpb_inst_0.INIT_RAM_22 = 256'hE528E7FFD4CDB7F30BA48007CD7FD2E3560FB5F80EC4BC8D7E7EA22ED9EFF3A0;
defparam sdpb_inst_0.INIT_RAM_23 = 256'hBCD00D396196BA4A616E37DC43E7BC736D1EA39BF83268ECCCE72E2E8C8BFE9C;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h85C90CB938BBC2386CBBE49C12157DEFC15DC1E246404A7A14D6AF44CC271BFA;
defparam sdpb_inst_0.INIT_RAM_25 = 256'hACC27066095CDC37D7C46C055D6DC7AC65223031B7A22B8C458E5B7DB842961A;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h24741E33C73663281298914A59DFF5C7B5A57F229E30B0BEAEA96A24F454A0CC;
defparam sdpb_inst_0.INIT_RAM_27 = 256'hB12FD41668C1603914F85A6519B1F276444C795B50EC0E352177DD18E1C2CA0A;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h887CE8557E6227820C648994F9E4C165E7EF7F6E699065CEF7B6C35AD9B7AA4D;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h1401AF1D339B0BBF0DBE4CC4C7EB050D7FA4ECCBC32400525BF6652099C790EF;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h06FAE3E39A703274DE974ABC7DEE0F7ABCD081938C9F5F1C16FCC44DB71E929E;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h7E89CCE423D055301F67273AE32A803D97BFFD731F970DBE16FF57E65DA0E721;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h68C14F975758A30F5E24C945EA3EA97055D773CC64B0D4B88BE9956408548DE5;
defparam sdpb_inst_0.INIT_RAM_2D = 256'hEFD15CF350C68CAE4D34471CAED7F9A232D819ABE012B7D71AE6EE81B86CA502;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h9B763A5F994939509DA7189D63460FBC037E58FFD47C7CCE6CA0C244454DCB97;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h6A1E01FC2CEC2D15ED24903AB40FC19EF00DB357BCC871E6CB658D61BE7A594A;
defparam sdpb_inst_0.INIT_RAM_30 = 256'hAE9EA482809A4A207D6846F6133F8067FBB0A7715FB0F8ACCC6C1C903F268267;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h5CF04DC0AC3E15449332C7AA92E6A82DA2C542F27CE682D621B62890698F188E;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h024B4F37260A2743B03F4E61BE0487136DDF037B3079EEB85969AFDCC002D12D;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h5162E21E811F761B5B0A8569996E6259D7B7DA74F6F7E5200A440B7A6215ED88;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h26C72E409C58727E83E0008A4F41EDFEACD8F13F16A313130164F13BF5C91FC4;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h285DFA2624BBAF9ABCEE15BFAAF9ADBFF09E150005A47FF2D40B90F7F7807CD8;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h637593FACF9FC4F3985193437FEB6763F7AE93BBD44AF5F764F0266F3DE582A6;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h0FE3B44CF50185300F7CDDFD2ED4712A9DBDD1BB2C0B24397DC633F6F1CA8A3F;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h191C5F566A348D0E004C1AFAE1EFE6FFF1FFF5B46CFC82B3FF4E3DC4FA8F8F8E;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h1DCD201E99EFDEDBEF40BE1F887ED57025CEFFD38D452F625906B5C98E2FF782;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h2706C417C16A2046F876D58A3B43BB2880E5DD72B7780D73156F4AA03AF23116;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h432609EF46E1EC6849D99571BEA008DE5F1C11F33E874BC74E08EDA98697F0C2;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h7A37381EA236C7B5AE1ECB8477FB80EF7BF22C79C0735144FAA80B4B386F7937;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h88151398A4312FBC0AB1813855E9081EFFFE4E4C7CA4DDCDDED4CCA1FF436157;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h81042198211F5A13D20D1916D03FCE023E58441E01F52B9CD2AD87FF2F70277E;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h7BD823B0DF8000D838264A49A897DC87765E1E0C3CFB79CF3E2E18A3EB473BE2;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b1;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'hA8FC435FC9DDCDCF9EABBC0003D527AF45757A5FCDF422AC06041980E7FEA3C6;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h3EA593012ED8AD97DCD8D82F9B42EDDAC4DAF2E3700F76C18439049A1FFFDC67;
defparam sdpb_inst_1.INIT_RAM_02 = 256'hD9E69F88F9A7BAFC6964C26D88E0624807C5340663867071C7FFD521B22CE3ED;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h5BBC88EC9ACA0925AEA4CF124989BF8E71A0FA01E3E7076D2FF922CA0B26F22F;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h9957A18FF51E96DBEA1C3CCBF4052CF8B215E827D2A3AB4D850CFC8FA4F53BF5;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h04F777C0717810192698B09330DC721BD7FB2F3C0CEB8EB4955BC9F84CCB6484;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h905FA7EBBF738642B20344A3FCE9AD717EE58B98102D077371CE03DDB1753B8C;
defparam sdpb_inst_1.INIT_RAM_07 = 256'hC362CFE7E91C441C19A8DD91ECA137129FD747B498FA9BD1F2853A1FCE9FC877;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h8C37E7C7681603BB1039A33CB0115B4489E20CFE0F71F9DB0DE66FDF9FF5D108;
defparam sdpb_inst_1.INIT_RAM_09 = 256'hD4678670E4672E9CAB00902A3F82BA3CD66E362A9C71B9040A765673F753839B;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h0D9AB54FFF0B9A3187009406799B2D06A1910D193FA87B1F25222818DC037A34;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h059C9D50FCE23B64BA802A0D204CDE9A7D1AED71AFE871D7EA172DFFBF856B8E;
defparam sdpb_inst_1.INIT_RAM_0C = 256'hA1D7A21B467783323ABC0208E9A3BBA103AAFDFAD4F15F221BC412BEFE607676;
defparam sdpb_inst_1.INIT_RAM_0D = 256'hB19F0D77D8067DB2EF9C4100120D7BA191266C0CF6B85F4E4CBDC6EAFFE3D26F;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h921EF623599CFC0510614AA1BFF3E94BD36246D2A6F3180BE13FF85714FF709E;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h5B75F67712B2A3C128AF9DFB502A973EB9BA40708D4A168DBF819FA85C77F5F5;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hB50DE7F77BFE571C09C80B5CB5BE754B80A30A9A2F44A46B01382FDDC5F186DF;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h5C28FDBA6BD885862F5058AFEFF7E5C8F82232001FE1CD9D9007C40C3011083E;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h4105E65FE349035C5DD58A7E4995A3FA4E539A04D8FB4FFCE8887EF08310EEAF;
defparam sdpb_inst_1.INIT_RAM_13 = 256'hBD30769ACB38695B71E1221C01A1AAB7E28F69CE12812099E4EF3171F21ABF7F;
defparam sdpb_inst_1.INIT_RAM_14 = 256'hEBAAC31B0A73FE741E9A722CB37E8F0B60948A5CDBB312C82538EE6FFCFDD83E;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h9B8F7575E682F03DE845DBB363E68775BA045AEAD7EFBEAC0E028F041E87CA2E;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h603B63CF56BEE8FAA0482672E6B790705FC00F556A70EF4AFB6A9FFDAA318C16;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h9D5D4BDE64AA0DBB202914DE3D9FCD11E26D0DEF3BB0CA4E9A1577F7392C8672;
defparam sdpb_inst_1.INIT_RAM_18 = 256'hF7CADFE77FB1DDFF716F528D5A19EFE3929FE25D3BAE55A6C1DC2157FB81DE39;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h3BF3C3FC8FCBE3FD000B48B5D302AE9E678744D44829E9FDCB4EC1A77FFE2278;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h1B564EE9FFEF7EBFFE25B869A7CD6CEB4035E87D7F66D2F7BA247E1F6E4777C0;
defparam sdpb_inst_1.INIT_RAM_1B = 256'hF33C13A50D7E5EA63285D902AB712581BEBBDE1B9FE26EFF7675EB0B8B5EA7FC;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hC7F87953F47F6ACB8100324E2B0C5551EE64F37821051683E408E06EB349103B;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h0078D870B3C32A6C618911C5241113A21F20F9E1E0C20E8026A09E952C0766A1;
defparam sdpb_inst_1.INIT_RAM_1E = 256'hE752C021B97329D2CB7A01DA656C1C17F022460EA2C175B17E0398C0225AFE4E;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h9BF4E7C81EAFEB5DFA9FD47092D97E2DD331E46AB359266D7BF1EF1D8885E7F0;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h7A43E215BBF489C56E554281424696710F98CC04F517DF98813D1F87090AD179;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h9774110B4B8BDF8207173DF580A0B27BF255E23944139DDD353B96F5E8E16EBD;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h33208FA834ABC8467ACD4CFBD1B73F6F161130218717EE7A618BBAA533783760;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h639031B21E56C50EE66D7075C1142EF3B67686E7E1AC4BD1CABF2DD7F06BE6A8;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h0CA17ED8A55756A9BB1668A8E83FFF98F098A4B815E945C036E31CE1946C500C;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h0B497EB332F49E5113364C62687F10386C2CB6AB36BA62825928525C962E88A6;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h0B684D7E1D5AFCE9C50E3233D98AC4408202BAECF7309BD263ED5E37DA8B4D2D;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h4787F71E7E6009818756DE5C2ED51622105783EF5DFFA5E2F57EB306AFFAFB8B;
defparam sdpb_inst_1.INIT_RAM_28 = 256'hB6669869F082464B5E12C4E2E130180F05062A4540B5FA091E5B522227476F18;
defparam sdpb_inst_1.INIT_RAM_29 = 256'hC51584D6282337327AC9472A546071E3A965A4540077EF80B6417EB6C9A1FC4E;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h234245DBFC1481EE45F8BD4FDCBBDC0678B586CE422F020762FAA1814DFE26F7;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h41A9C9E7B7870E16B6BC41654CE3918F1164FCF2C2EB96EB4E2B6EC83CA2ECD1;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h033F75FCB3713024D390926DB27659E3A15677FFBA5EE6326CC871FFC5AF7409;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h0E10C84AB134BA75CEA214819B85C97F20E3E66650FCD54F6B7C98F10A0AC6CE;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h3C13728B08DB96304B5AED0DF9B772D1F2F9FEA2020140E761C5EDDCDE2B7F98;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h7855F7032A3EDC640751F4F90A43714F6E49E8C04989C031BCE6BAAF49983F2D;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h7245DC7DFEC6779980028450223BDA6E56EBB0103B3E9C767DB02656CEA12481;
defparam sdpb_inst_1.INIT_RAM_31 = 256'hE009400632D3CC74056314D46DCD208E73D70E07FC77FE7AC8260D3073ED4988;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h083C7EFBB0F5E287929D15E8054068E1B8CB6DA7907B340B7944EFC1696875E3;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h89F19D1AE11AF2DC7435C4A5A4F4F8F1D98CE0F266F9BC062911A8DE045B910F;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h3718DC619B0A8944299CE59FD24AB2AB2EB3572538B66C80450C98EF61D4C50B;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hF92ACBB820F3F62019CC5011EE0D3EEAFDA7772218501991BB073A1639950A93;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h6220346F572B13B0B8F12506BF7EB82AB637AF6709C86A9F6597CB20533C8D28;
defparam sdpb_inst_1.INIT_RAM_37 = 256'hFF98F8B2F9D0BA515A5B8A88F1ACCFFF2AEC4F902B7250CA30357D78852DD255;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h3DD23C8B39D4C58A15DA3C01D8EB174A52CD49EDE1701E4AC93248BCD38F80DC;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h8DE5CD9C84E07E61DB87513B5E5D803EF483106313C1360CE4D8E406C1479022;
defparam sdpb_inst_1.INIT_RAM_3A = 256'hD04596F7850930310E68A97DAA7AE3DF5A39BA3A2AFB6A0E3231E53B1EF8A4E8;
defparam sdpb_inst_1.INIT_RAM_3B = 256'hB8E99247D28E08F36313E1510F46785D89E981972786EEE15195E7CF38D50702;
defparam sdpb_inst_1.INIT_RAM_3C = 256'hEF4D9FC98A29DAE985778682A97FEBFD7DBEBC385146E56C780BA2E1486675C5;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h1224BE97071409E38F338D22400D7FA15065864E97A450A7F6D8CCF0EE4DE2F6;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h622E2A1D593D3F8A4A6CF7BBC0EC3EC84EAC75F4B1830D484E4ABD7ACFCC0B1C;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h695CA48B1B2B7D6931CB8A2347DAF8D493AA4015C8235630852C519897182E3C;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b1;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'h97D3583046BFF483FF20100138801BFFFFFFFFFFFF7FFDFDFF44021ABFFFE146;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h166B114806197B011FE2000A7DEC09AFFFFFFDFFFFFF6FE3AFEF10080E4BB2D6;
defparam sdpb_inst_2.INIT_RAM_02 = 256'h68D788400013F7800FFD000769FFF002BF7BFFFF7B860C03C5DFFF0200C7FFFC;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h4F877F000102FEE801FA0800F7DFFB80637EFFFA82028004861CFB62880184F7;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h2F7C3E060441BD78414F840037DD7FFC4010F05C9000040011C4407D6E6048C9;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h012936F322027AF6224BFE0003C767FF4100772B00B200020115401FFFEFDC00;
defparam sdpb_inst_2.INIT_RAM_06 = 256'h00259D1E201246BFE007E7000084E0BBB800473A1864000020003806EFCB70C0;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h80001218800C522DEFC41EF8206000AFE0040DBF9A0600000000906E5A677F88;
defparam sdpb_inst_2.INIT_RAM_08 = 256'hF4B48B80C830040DFBF829FE80106AA4FD001C17FA50000055280100777FF9FF;
defparam sdpb_inst_2.INIT_RAM_09 = 256'hBED27C052D0033C02D1C004BFC03FDA43FE9FEE9FF7B06004000C00800BD7FFF;
defparam sdpb_inst_2.INIT_RAM_0A = 256'hFF7FF4111182118CEBB8E60F7E401FCF2DBF3F7F977FB480540B0030417BF6FB;
defparam sdpb_inst_2.INIT_RAM_0B = 256'hEFFFFB5C96124483FF3F7C405FE820FFEB8FDB67FFFFFF80000023500C2FEDAF;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h70FEFF8EA241280817BBF7D4017F23E5C60E185DDF7FFDF0000000B500006CED;
defparam sdpb_inst_2.INIT_RAM_0D = 256'hEFFEFFBFEFD434C30BEF7FF988175C533BCC39C27FFBDFFE000078100081046F;
defparam sdpb_inst_2.INIT_RAM_0E = 256'h6FDFFEFFEF6CC480CA4733FC080DFFEBF4BF2286871AF6FFE0102F0C28E8884F;
defparam sdpb_inst_2.INIT_RAM_0F = 256'hA7DBFF3FFFFFB9804832CD2EF8427EA9F3559E3AF98780BAFA100ED13000B023;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h00CE1AF29FFFD3D480CBFD7FF00801FFDDDE17BED7B4CC01FF08E26AB9000100;
defparam sdpb_inst_2.INIT_RAM_11 = 256'h00077FFFFBFFFDBF5A904BBBCB810813F279E727FDC1F2C003F4600D0D9A0010;
defparam sdpb_inst_2.INIT_RAM_12 = 256'hA8000A7FF7EFEF7DF20268DFFF7CC2115F1E39E8116586EFE40F208E01333140;
defparam sdpb_inst_2.INIT_RAM_13 = 256'h5C800003BFDBFF97FFF48F85F7DB00002F6D309734EE85FD7F02F00695EAA695;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h649988017EFFDFF7FEFB005B7DFFF80000FB09209481314B603C1D842CE5EF9D;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h723D1F00003F6DFEFFFFD2867DF38714010DF1E197FB226A6481F8F000DB93E4;
defparam sdpb_inst_2.INIT_RAM_16 = 256'hE85863048C17BFFE3C9FF7D505FFF780C4085F8609327D7AC993879F80079148;
defparam sdpb_inst_2.INIT_RAM_17 = 256'hB3D1028000DFBFFFF77DF7F903FBFFF6400E0FC0CD4B47F2038086197E0170ED;
defparam sdpb_inst_2.INIT_RAM_18 = 256'hDF136604000007FBC7B38FF6D5033B74600008483A5B64733D0DF73B1F740F78;
defparam sdpb_inst_2.INIT_RAM_19 = 256'h9726E5B022801C53EF66E557FD0FDFFFD1001000833205CBD511DA9DB1FEFFE4;
defparam sdpb_inst_2.INIT_RAM_1A = 256'h50AE844E41400141FF7DE375FBC75FFFFE88080600346584942013AB59C3FFF6;
defparam sdpb_inst_2.INIT_RAM_1B = 256'h56856097B4004100FBFDEC3AAFC6EBC9FC880800130EA4610E7680910E98221E;
defparam sdpb_inst_2.INIT_RAM_1C = 256'h19EAFB1B9C6231021FF7FFE776FE6A66FFDF0B640001A535EAB8DD90B2A9E089;
defparam sdpb_inst_2.INIT_RAM_1D = 256'h584671771185830000FFFBFF18FBFCEFFFFF920E63001E38554FF1F632E97F37;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h0E70A423C72CEC08002BBBFFF37DDDE5B887BFBAFE9020E7E44E281F339DD0E6;
defparam sdpb_inst_2.INIT_RAM_1F = 256'h0E1CD1DE12F7AD30300279FFF80B16FA237A77DFFFF38018BBE8F7CDF375C71D;
defparam sdpb_inst_2.INIT_RAM_20 = 256'h0024E1925D51C8B9A0100FF7BBC4B9FFE06F37FFDEE6301798F76725F5CB19B8;
defparam sdpb_inst_2.INIT_RAM_21 = 256'h7001ECFDFBED07473268416FFFBD2D36F833FFFFF7D1BE1491545ADC3F0033FB;
defparam sdpb_inst_2.INIT_RAM_22 = 256'h230A32D7EA60331E127C800FCFFFFAA7FBF05F9DFFCD38B1AF96E7C1BF738D09;
defparam sdpb_inst_2.INIT_RAM_23 = 256'hFFB04878E1C6F508D98243D4FFEFBE3B6FB11CF3E2CCF0E73D5BA70E4AFA161E;
defparam sdpb_inst_2.INIT_RAM_24 = 256'hD50B08D31942A63916953DFD3FFFFFEFC17FE43DFFFFABC97ED334F3AF5699B9;
defparam sdpb_inst_2.INIT_RAM_25 = 256'h9DACD9A5932A1E2ED5765B0CBD6FE7ACA413FE00FB9FF4329E7FA2622EA51E1C;
defparam sdpb_inst_2.INIT_RAM_26 = 256'h4BFDF1F989B59C6090D7E825947FF5FFBDA5FFE36FFF9F42650804494CFD5C3A;
defparam sdpb_inst_2.INIT_RAM_27 = 256'hE08C268F814B0FC5D70ED89E07B7FAF7D64C7DF90E7F75DC8B747219A601B1DF;
defparam sdpb_inst_2.INIT_RAM_28 = 256'hBE7284ACFF42107D4973EE05001F7FFDFFEF7F6F9C6FDDF1356ADFAB75B01A8D;
defparam sdpb_inst_2.INIT_RAM_29 = 256'h60373AA88FDE6580E239B1B2C81070FF7FE4ECCFFD03FFEDA42259C22CB1602C;
defparam sdpb_inst_2.INIT_RAM_2A = 256'h056FD31749FD51E90093576DB8000D957FDC81939F7900E7E9021661B1B563A3;
defparam sdpb_inst_2.INIT_RAM_2B = 256'h81714AE689B86F148013B7F5E9910020AFBFFD771FF98401680000D42EF5DDE3;
defparam sdpb_inst_2.INIT_RAM_2C = 256'hEB66E5C810B3E2BB560632657D980031DC3FF3CC44B31CC774160030F7572934;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h07A7C1F84A527C3107F4D596774BC0220C41FBABE012B9C1A50900019DE32833;
defparam sdpb_inst_2.INIT_RAM_2E = 256'h8508383A3BDB474401B4945533D7F60002FA2FFFF43C6F1E20562444406E9818;
defparam sdpb_inst_2.INIT_RAM_2F = 256'h1A4606FA845FECF40BC236874F115430003A74F7BEC851F9C89A2001BF80B423;
defparam sdpb_inst_2.INIT_RAM_30 = 256'h15D593375F56D998025526DD34E1B983801FC10FDFB0E8AF1E40C0403EC495A3;
defparam sdpb_inst_2.INIT_RAM_31 = 256'hE900A396D195333390CAFE9844894C5FBE06B7D1BFEE82D77C9054002FF1E6D8;
defparam sdpb_inst_2.INIT_RAM_32 = 256'h9A4B0AA0257110C750001E79FE467C43877FFAED0FF9EEB85FBF0008803D593C;
defparam sdpb_inst_2.INIT_RAM_33 = 256'h378FF0597FFAD9B8C7037A1F36A8DFE3ABBFE3AC91F7FDE003D9C80020160E52;
defparam sdpb_inst_2.INIT_RAM_34 = 256'h9740673B7CC7CA81F0407FF3BB40A3FF219A879DC59FF313007F8F00000979E2;
defparam sdpb_inst_2.INIT_RAM_35 = 256'hC3F53F8E6C47A05AFC1E0AFFCE0F7C7FF99780BD48D5FFF2D40BF96080407B1C;
defparam sdpb_inst_2.INIT_RAM_36 = 256'h8DB2A68D758FC30C100F90BDFF0EC91FF7CEF202C2FD8FF766F0379D000103D8;
defparam sdpb_inst_2.INIT_RAM_37 = 256'h78CA42E990A580CFE083FC02FED781617DFECC0E6479B5FDFDC6BBE8F000227F;
defparam sdpb_inst_2.INIT_RAM_38 = 256'h1A6A8F74AC2449F7FFBFDA811FEFE7FC0FFFC7903F6C788FFF6E0FC70E901B0E;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h1FF23687554EA687FFFFFE097FAED550003EFF1511156F399FE6B6C9F1A80022;
defparam sdpb_inst_2.INIT_RAM_3A = 256'h0324B1964F637FA1FCF7DD80C4BFFB80002F3D7CD53F87A60E7F4EA01F0E0080;
defparam sdpb_inst_2.INIT_RAM_3B = 256'h2325FA0D1302BA2739D99971051FFEDC5F0D5CFBC7722EA6D2E8FDBB86B1B404;
defparam sdpb_inst_2.INIT_RAM_3C = 256'h80135F60B34FD350591ACB8440007FEF7FF2C92FFFB863370C454FCB386D9728;
defparam sdpb_inst_2.INIT_RAM_3D = 256'h0C0433FF40C7CEC912B001380202FFFEFFF94181FFFB9E4CCE7B2FEFFF0BCCB0;
defparam sdpb_inst_2.INIT_RAM_3E = 256'h3104219FFFE39D0B06AB12169000317DFFF6484EBFFFD41DE84F39FFBF722792;
defparam sdpb_inst_2.INIT_RAM_3F = 256'h8FB823B6E7FF831D033C3A0993900108898D792BF37FE6F0314E0B5B7B673BFD;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b1;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'hD9BC00DFDFDF7E0C5AA2CB800B33000001C7BC0FCC0BDD57F87A7396F7FFE377;
defparam sdpb_inst_3.INIT_RAM_01 = 256'h2F1F83012ED9A5FAE249A29E2E06F4000505579FF000893F7FC33766E3FFDC67;
defparam sdpb_inst_3.INIT_RAM_02 = 256'hD9F9BF88EFCFBAFE91590D3B80E0E20006BECBFFB980867E3FE41202B7FBFFFD;
defparam sdpb_inst_3.INIT_RAM_03 = 256'hDBBF06CC92DA0925F93446A3398B3F8E71F2B9FE7C09E3E398FFDCA0F47DFFCF;
defparam sdpb_inst_3.INIT_RAM_04 = 256'h7BD7F87F051096DBE7E17C3D3385E4F8326FB8000229CF7E79DFFF713118AFFB;
defparam sdpb_inst_3.INIT_RAM_05 = 256'hFEF77F0E7178101836FF251F9E3C721FC7E031200C39B2961BC5FFFF96FD6F7F;
defparam sdpb_inst_3.INIT_RAM_06 = 256'hCFFFA6F05F230642920FF630A8A7AD81FF79ED981E34EF085F2F3FFFFEF67DB3;
defparam sdpb_inst_3.INIT_RAM_07 = 256'hF29FDFFE1790540C1920DE3072ACF7191F8E3D749E46B82EDC5615DFF7E7BB3C;
defparam sdpb_inst_3.INIT_RAM_08 = 256'hAC907FD7D0F6001B1039A3C5B69EC744C1F2929E0E5B1825EEC155C99FFF19F7;
defparam sdpb_inst_3.INIT_RAM_09 = 256'h0FCE9BF3FF2D2204EE0040F46921D9FCD58DC6D6DFA19803FE49B0DCBFDFFD80;
defparam sdpb_inst_3.INIT_RAM_0A = 256'h9FC8AC3FFFF2F8018700000792AC5B3EA5A91A487FC23700FE30881B498B7FC6;
defparam sdpb_inst_3.INIT_RAM_0B = 256'hF8BD671BDFFFE700BA80A20F353A3545FD1F944C9FF05FD407E6640045EC7FF1;
defparam sdpb_inst_3.INIT_RAM_0C = 256'hFE1D2C783FF7F8F2009C0200FA3C9C84EFBAF70013FD44A2003AB480018E637F;
defparam sdpb_inst_3.INIT_RAM_0D = 256'h4E605DD5F3FD764ECFACC10017FFB7E88FFE7FF0FA7FBF3E40001299001C7CFF;
defparam sdpb_inst_3.INIT_RAM_0E = 256'h67E100C5CD43FFF8F0714EE537FDAF0F909FFEFD6C4FED57E100017B0000CD40;
defparam sdpb_inst_3.INIT_RAM_0F = 256'h5E0A086DEDFC1C0E37A09D7B502FFDC1C385FBDFE9B9FA43FF8020333C000A00;
defparam sdpb_inst_3.INIT_RAM_10 = 256'h07481007A76E826FF0380B5FF5BFF80412E4F4FFD12A5AF0FF3806062BF00120;
defparam sdpb_inst_3.INIT_RAM_11 = 256'h002FA0427B46F341D04FDCEF7FF7C26FC0160DFFF82B22506FFFC0003A310800;
defparam sdpb_inst_3.INIT_RAM_12 = 256'h41029A00236F4F8E0261637ED797FF8ADD1994FB2700B705877FFF90453BEEAD;
defparam sdpb_inst_3.INIT_RAM_13 = 256'hFD3066B0013BDE43401824EF73BFFF417CDCC423ED7C8A01B212CD7042DC5F7F;
defparam sdpb_inst_3.INIT_RAM_14 = 256'hFF9AC3C28073FE8CA581D25EFFFFDFF46B45C3C3240CDE78392011DFFCFF59FF;
defparam sdpb_inst_3.INIT_RAM_15 = 256'hFFFE7C793682F38A41B0E43957FF79FECF8CF398201043690F9400FBFF87FC2F;
defparam sdpb_inst_3.INIT_RAM_16 = 256'h8EDF63CFB6A2FEF4C2FD90421CF7FFEAF2514504C00600455BA9C002FFF18AEC;
defparam sdpb_inst_3.INIT_RAM_17 = 256'h52BD6BDE69EE0DBFE0C369C232FFCFFE0DD3F5C39A99308C6E5D348007FFE465;
defparam sdpb_inst_3.INIT_RAM_18 = 256'hFF17D7E77F879DFFFE05AC7D0A7FFFFD6D1DA351D981222AB13F0DC0007FFE2B;
defparam sdpb_inst_3.INIT_RAM_19 = 256'hFBA0BFFDCFC36FFFFFF37F737321FEFFB887F231AAB800004586E1CE0041DFF8;
defparam sdpb_inst_3.INIT_RAM_1A = 256'hFF57DE69FFEF0D7FF7DA20432BDF9FFFBE86FF47D141C0003317F85AE802883F;
defparam sdpb_inst_3.INIT_RAM_1B = 256'h0CFC20430D7E6BEF7FFA21A5D5DDA2EDBF438C5CFC001E00026BBFB7DB420003;
defparam sdpb_inst_3.INIT_RAM_1C = 256'h00079DDC3C7B76145FFFC401DD9E172FFFD9E43F724F6180600EEBF74CC91004;
defparam sdpb_inst_3.INIT_RAM_1D = 256'h000607FA8B3FF538FFF2CC01511605C1FFFF0D13E465F7180680C5BEBBBF66A0;
defparam sdpb_inst_3.INIT_RAM_1E = 256'hE750C01F2A921519860DF620070742E90FFFFAAC0143F640FE0395A7CDE9FE4E;
defparam sdpb_inst_3.INIT_RAM_1F = 256'h1BFEF7C81F70F4AE92E028080AEC142618DFFBFB46DC522447F9EF9B75489FF0;
defparam sdpb_inst_3.INIT_RAM_20 = 256'hFAFFDFEA4408C67D959C25404047238AF147FFE7A0C8231AE4FD1FBCC6A612F9;
defparam sdpb_inst_3.INIT_RAM_21 = 256'h7FFFFEE0DE3848511BE9020080A0FD9697DC7FDC6D358C01CEC7F7FF0607E58F;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h0DDFF04038DA707D5098BC0241B57F9981C70FDE6D1E102D8B7E4FEFC6206853;
defparam sdpb_inst_3.INIT_RAM_23 = 256'h902FDE003C95A7C4FA9B0FF1010C7EF879D1F81D05F3620DDA7D62FFCEF40B31;
defparam sdpb_inst_3.INIT_RAM_24 = 256'hAB820020BA65AA3EF709411E403FE7FBE0756A87E83296BBC7E2121FFF834137;
defparam sdpb_inst_3.INIT_RAM_25 = 256'h65B80404B31958DB771E3C1DD87DFFFFFF864E19C903175EB0601ABB79C0F0F4;
defparam sdpb_inst_3.INIT_RAM_26 = 256'hED8BC00101B353B272F771F0068FFFFF7DFF45F2C080D3C3B80250C325741EAE;
defparam sdpb_inst_3.INIT_RAM_27 = 256'hF8DE8600007E2F724D66BB22012DBFFDEFEFEE2BEC003BAC91A79127F805004B;
defparam sdpb_inst_3.INIT_RAM_28 = 256'h878E2BE80003AD14EDFCC45C1E0FFFF6FBF9FDB045B80AFBE2BB2B145F199038;
defparam sdpb_inst_3.INIT_RAM_29 = 256'h6ABBDA86002239AF3715846C33F00FFD56DA1BFBFC2FA79611DE5D9E1B600007;
defparam sdpb_inst_3.INIT_RAM_2A = 256'h0C8D8608F610AE75F1C76AA21486C2F567626025BBFCE3FD5C31381B21B60000;
defparam sdpb_inst_3.INIT_RAM_2B = 256'hC1DC110E8F871FE49DAE7A3221EC6F80FE9901083C0018FD6329C18647B4F400;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h03366278A8B136F9DFA2794BAEA0F61B0EA100004120065B025095E022856E00;
defparam sdpb_inst_3.INIT_RAM_2D = 256'h86931A0BDA8BBBFC23D50744392234C0E034002000234B45ADABEECBDDD8AD6E;
defparam sdpb_inst_3.INIT_RAM_2E = 256'hCF17626AE2B07EF78EB42A651FBC28CD0FF800200201022611327FF3DEFF32A7;
defparam sdpb_inst_3.INIT_RAM_2F = 256'h47FBFC95FCC6C79BF865C4590005394939BEE88009844021E63DCC1C9586EBD8;
defparam sdpb_inst_3.INIT_RAM_30 = 256'h41BEF994521BAF3FFF0C98AE7CB68A4255244C107B3EB4F63F373A814A083104;
defparam sdpb_inst_3.INIT_RAM_31 = 256'h23061FFB592241F3FE83DA5A795A004D565E01F7FDF7FF7AE9E6DCAC1FAD01C3;
defparam sdpb_inst_3.INIT_RAM_32 = 256'hBEB9010020D263DF2D00595F3FBC130CCEB34C84EF85FFF9FEBA923C9FC77463;
defparam sdpb_inst_3.INIT_RAM_33 = 256'h1B5B80A80221053CF0E807142BB5740F6C84548A6400CFF93EFE0B69CCE0AD07;
defparam sdpb_inst_3.INIT_RAM_34 = 256'h0CA5F80223EB9901E78201A3441AE28CEC3B8A20EF81B07FBEF749BCCD2B3480;
defparam sdpb_inst_3.INIT_RAM_35 = 256'h27FBEBB800FD297BE43C101E3446B0D2C9FA867FEE20025040C8CA0C1B8EF17C;
defparam sdpb_inst_3.INIT_RAM_36 = 256'hCCFDCF1F572FD11709772907C2D7BF4FA736E61F6849FE8262204101A4B5FAD7;
defparam sdpb_inst_3.INIT_RAM_37 = 256'hFF99DC71FBD7E3CCE0E67E88FE37AACE581A5756CE85DB2A000802D08E5B6FF7;
defparam sdpb_inst_3.INIT_RAM_38 = 256'h07D3565D4BFFFA1ECE8EE7B5DF03A69E3F1BCB3512A38895C03A004CD7EDE468;
defparam sdpb_inst_3.INIT_RAM_39 = 256'h791938EC63F7FD8766040C1FEFE23AD7251AB17754E705420AD0E00281F463EE;
defparam sdpb_inst_3.INIT_RAM_3A = 256'hF2C86EB6C33FCFC1FB213AE277FD030C51158C8422E2A976085DE5BA7EE7C64A;
defparam sdpb_inst_3.INIT_RAM_3B = 256'h6207B18998C1F70C7AF3EE7570B9807974B115FF7CAE5B719B917FFF7FFFFB2D;
defparam sdpb_inst_3.INIT_RAM_3C = 256'h72CD82F32CF02D80000D941966801C01B532FA5AE1A1AAAF924CC5BA4BFE7AA4;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h9785F81845BCA4010FDD60332C000020FEA9E7BB27EEA97F5401CFCF03FA8510;
defparam sdpb_inst_3.INIT_RAM_3E = 256'h24B9F0197B7E68000BF1C5BD3A4C0A404FC917922A15C6D83897B71A303BF420;
defparam sdpb_inst_3.INIT_RAM_3F = 256'h000FC6CF7148EB0931DC09001727F88093FC6A00EA09B1170888C25FA0E17040;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[29:0],sdpb_inst_4_dout[1:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[15],ada[14],ada[13]}),
    .BLKSELB({adb[15],adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_4.READ_MODE = 1'b1;
defparam sdpb_inst_4.BIT_WIDTH_0 = 2;
defparam sdpb_inst_4.BIT_WIDTH_1 = 2;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'hFF3FFE8D656E1F1CE2B2EA0128D05BDF8C657F35344B780535EC15808444041C;
defparam sdpb_inst_4.INIT_RAM_01 = 256'h8C33FF0CFCC66FCD5181E2AFA4D99F31133F3FFB9428350AD493363BABFFCFF3;
defparam sdpb_inst_4.INIT_RAM_02 = 256'hFFFEF29AAE664D81105CD11EA2A2949471A30780D91B04355B151707C5DCC834;
defparam sdpb_inst_4.INIT_RAM_03 = 256'h33DF7BB5BCC27483A5EB741D173D737B1733B3BAA950CE224D47DA4F9B27BBF3;
defparam sdpb_inst_4.INIT_RAM_04 = 256'hBECCEEEBAE6A8950F09002F9C97A8FD8FC35FE91484CD897FD3C3FBBB8B05F0C;
defparam sdpb_inst_4.INIT_RAM_05 = 256'h79F832A663E7172550FD9180DB30AC5B2FEF34F7EDAEAAC1985682E19A692BA6;
defparam sdpb_inst_4.INIT_RAM_06 = 256'h9CAF6EAAEB69596920D50588A5BB5F2423862F6822401063DC588F426B0EF82B;
defparam sdpb_inst_4.INIT_RAM_07 = 256'h1BB6B1AA72CBFE545001335B34EAA5B0DBACBFBCAA0A64841D459221541BDD5A;
defparam sdpb_inst_4.INIT_RAM_08 = 256'hDB1A6AA5961956955457FD1E48DA8ED8695379A1DB5F94DDE38CE29C13BE36EB;
defparam sdpb_inst_4.INIT_RAM_09 = 256'h1F7B7DEDA63A83959034194FF989B4134A9BEAFB5AE2A59433D31DAD659A23E1;
defparam sdpb_inst_4.INIT_RAM_0A = 256'hEDE7191459429906A51110FAABF922B3AAF508223D1E8BCA1DC366C31EF5F29F;
defparam sdpb_inst_4.INIT_RAM_0B = 256'h5A5F7AAA45691891611C420BF3FDA6AA3066A4BD166514451833E5C3D8E6C2D8;
defparam sdpb_inst_4.INIT_RAM_0C = 256'h6AF0534205010441411151D8C8E6CF93908FC6D98F74097F940288FBD8F65071;
defparam sdpb_inst_4.INIT_RAM_0D = 256'h1F04551A6F0D80D86FC80F0CD5C0E2C9A567996B09A40E354100FFAA7AD80E6D;
defparam sdpb_inst_4.INIT_RAM_0E = 256'hA996BCF00403C01500CF15C4F70F36002C8B82D4682772F8DCD9533D981C6908;
defparam sdpb_inst_4.INIT_RAM_0F = 256'h6B5BF41544555B404400100CE1F83E489AD696A61A5050D47FCD12F7D940040F;
defparam sdpb_inst_4.INIT_RAM_10 = 256'h52D6F1AFF0F07503C08FCC30031000FF9A8CF4DF471C13128FF3BE0B1862517A;
defparam sdpb_inst_4.INIT_RAM_11 = 256'h4A3A9480104448D003F06F32CE2FCFF76AEB95D425A177DC3FFFCFCAFBD55054;
defparam sdpb_inst_4.INIT_RAM_12 = 256'hA817FBF6DBAFEAC3C03FF3C03CF08F12FFECCE94A1176BB537EBED76D80D35D8;
defparam sdpb_inst_4.INIT_RAM_13 = 256'h71F83AE6BDD3040510C3FB88B99998ADBEE19A91599591104BEFEEE9AA239198;
defparam sdpb_inst_4.INIT_RAM_14 = 256'h1151559141A6AD19AA6EBADBEFEEBFB3BE38FCFBEA3DDBD8CC06FE02F421C486;
defparam sdpb_inst_4.INIT_RAM_15 = 256'h2E96D9F4FCFFF14307C333FFAEBBB4114A64A5605561D00C29BEE7F652A6A156;
defparam sdpb_inst_4.INIT_RAM_16 = 256'h514E5004405599A5A6965EF96E58A9EBC33E9F30F03F64E606D498E2C4547308;
defparam sdpb_inst_4.INIT_RAM_17 = 256'hA73530E72BE47E0EF3FFEAC4B68298E9991155468559D41103FEF69A64194956;
defparam sdpb_inst_4.INIT_RAM_18 = 256'h851640554401B45625591DF16413105AAADAD9EA0307C3E95EEE900E4AF13848;
defparam sdpb_inst_4.INIT_RAM_19 = 256'h78F559F121AFED6AB2ACBCFB2691D5E550444C185044C717003CB8255C015504;
defparam sdpb_inst_4.INIT_RAM_1A = 256'hD7008D0F0C3F0144635343904911003405467B8A67AF001C3CE4DC6DF90666A4;
defparam sdpb_inst_4.INIT_RAM_1B = 256'hFAEAB3F32F30B1715ABB9A1B95A14D4551400FBB05FF0FC10B233EA1351FCE03;
defparam sdpb_inst_4.INIT_RAM_1C = 256'hCFCA8CFBFFFFF004F0CCE0F01010F03F200010096E67A030151D329D834DB702;
defparam sdpb_inst_4.INIT_RAM_1D = 256'h40E8D852558B78226C0AA96B79490E613B100EE22FF2FF3FEF8BBEBA0103D8C2;
defparam sdpb_inst_4.INIT_RAM_1E = 256'hF2ABBF9BE9FAEABC07E1C4F8CFC0FC0EE8C2333C04656AECCC01540FD4724D11;
defparam sdpb_inst_4.INIT_RAM_1F = 256'h96FBA62A148D9C408FB316AA56AB4520FFCBAEFD99EABEAEAAFB25DA992F0B5B;
defparam sdpb_inst_4.INIT_RAM_20 = 256'hDA8955965996AAA7A2BBAEFEFF6AEA6AAAAEAAF98BF33415AA03014981CE360A;
defparam sdpb_inst_4.INIT_RAM_21 = 256'h3C931B0CE63720082BEC601545282854B0B6AAABB95A95927AA92E6A9AA26FDA;
defparam sdpb_inst_4.INIT_RAM_22 = 256'h955C5145D866AA9A5AA9696A9AAB646AAA55556556AE9FF3116988C2596A53D2;
defparam sdpb_inst_4.INIT_RAM_23 = 256'h3836B01F6B62F2EDFEF1D97C90000F00430DB9658AA0012621D24549645416A9;
defparam sdpb_inst_4.INIT_RAM_24 = 256'h555F1A5C5C0C08151162112D8158440568410D017A55598FCBCC1DACC5A656A1;
defparam sdpb_inst_4.INIT_RAM_25 = 256'hA903C11C5917362AC3C57490F0113561F50F0FAE4C91145D1CC75345300843FB;
defparam sdpb_inst_4.INIT_RAM_26 = 256'hFAA4C47302CC3FEB1E03D11004430410D30C0C3C0CCE0005575AF001BBC11ABA;
defparam sdpb_inst_4.INIT_RAM_27 = 256'hAAA860FADC75000727117BC11EBF0C0C37E730482239B0C0FF9FEC7C0F3F040F;
defparam sdpb_inst_4.INIT_RAM_28 = 256'h2E515FEFB76A6F8BCBA3F0F3030F83CB8EF03FFF3BF3A383C3F09AE405A68366;
defparam sdpb_inst_4.INIT_RAM_29 = 256'h555DBAA40D4E0B0DFE8205B12F4230D00DFF7FC8E8D3EDEEF6E5EAAFBBEBA8BF;
defparam sdpb_inst_4.INIT_RAM_2A = 256'hA665CDF2CA6EEBAA0BA5E6E9CFFCFBBBFBAEFFA6BBB62EADABF0BF016AC056A8;
defparam sdpb_inst_4.INIT_RAM_2B = 256'hAAF1652F9A93F9E5D5AF60641D6514F00C0FCA6666D92CAEAAB6769A1A669A1A;
defparam sdpb_inst_4.INIT_RAM_2C = 256'h100EE43F9A791D656C065A5554DAFA666FAA9A58226B665A1568BA5DAC1AEFD5;
defparam sdpb_inst_4.INIT_RAM_2D = 256'hB142EC15A6BA68CE93A20F30DF43F2DB802EF3FE9259A1CDC8245AAA60450101;
defparam sdpb_inst_4.INIT_RAM_2E = 256'h000DCF32756543F8C4014CC01150501460565545348515FC745F8C165578C54B;
defparam sdpb_inst_4.INIT_RAM_2F = 256'h1BB0857F4707AA75510D3ED33BA2102C64C3F33EA5594A53229962010C43036F;
defparam sdpb_inst_4.INIT_RAM_30 = 256'h3A2AF0BA6563DF23FCFE83A0CDF0173305C00014F2FD5EF7CBFFE9C3BC896EA8;
defparam sdpb_inst_4.INIT_RAM_31 = 256'h9A3C5BB046AC129A6A4440BFDDA57429B1A3C2199BAAA8018E775A28C1FBCFC0;
defparam sdpb_inst_4.INIT_RAM_32 = 256'hB925A564993FC61A668E5E6096A66EF7217B3FBFB8FFFFCAFFAAAA5DB8AD9210;
defparam sdpb_inst_4.INIT_RAM_33 = 256'h00000000000000000000000000000000000000000000000000000002B7803FAF;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b1;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'hCFF3583040000B7FFF20100000001BFFFFFFFFFFFF7FFDFDFFFFFDE54000017A;
defparam sdpb_inst_5.INIT_RAM_01 = 256'h1DFF1140020004FFFFE20010000009AFFFFFFFFFFFFF6FE3AFFFFFF7F1844007;
defparam sdpb_inst_5.INIT_RAM_02 = 256'h80FF88400000007FFFFD000290000002BF7FFFFF7B860C03C5DFFFFFFF380000;
defparam sdpb_inst_5.INIT_RAM_03 = 256'hA0077F0000000117FFFA0800C0400000637EFFFA82028004861CFB7FFFFE7B00;
defparam sdpb_inst_5.INIT_RAM_04 = 256'hD0803E0600000287FFFF8400202200004010F05C9000000011C4407FFFFFF736;
defparam sdpb_inst_5.INIT_RAM_05 = 256'hFED6C6F200000009DFFFFE0001382B000100772B00B200000115401FFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_06 = 256'hFFDA621E001000001FFFEF00001314480000473A1864000000003806EFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_07 = 256'hFFFFEDE080000000103FFFF8206F6EE070040DBF9A0600000000906E5A7FFFFF;
defparam sdpb_inst_5.INIT_RAM_08 = 256'hFFEFF47F080000000407FFFE800301EA03801C17FA50000000000100777FFFFF;
defparam sdpb_inst_5.INIT_RAM_09 = 256'hFFFFFFFBF100120000E3FFFFFC030074C015FEE9FF7B06004000800800BDFFFF;
defparam sdpb_inst_5.INIT_RAM_0A = 256'hFFFFFFFEEE401010444719FFFE402034224273FFB77FB480540B0000417BF6FB;
defparam sdpb_inst_5.INIT_RAM_0B = 256'hFFFFFFFFFFFC0000000083BFFFE82001502044AFFFFFFF8000002350002FEDAF;
defparam sdpb_inst_5.INIT_RAM_0C = 256'h71FE7F9FFFFFC8000000082BFFFF237427F1D4A0FFFFFDF0000000B500006EED;
defparam sdpb_inst_5.INIT_RAM_0D = 256'hEFFFFFFFFFFFFE00000800067FFF5C204837463D81FFFFFE00007C100081046F;
defparam sdpb_inst_5.INIT_RAM_0E = 256'h6FDFFFFFFFFFFFE008000803F7FFFFE00336FFA3F83FFFFFE010340C28E8004F;
defparam sdpb_inst_5.INIT_RAM_0F = 256'hA7DBFF3FFFFFFFFE0800000107BFFFAC008DFFF617677FFFFA00090FF000B023;
defparam sdpb_inst_5.INIT_RAM_10 = 256'h00CE1EF29FFFFBFFE00000000FF7FEFF20033FEEFE6833FFFF00028EA3000100;
defparam sdpb_inst_5.INIT_RAM_11 = 256'h00077FFFFBFFFDFFFE000000347EF7FFFA87CB672BE20C3FFFF44010D7720000;
defparam sdpb_inst_5.INIT_RAM_12 = 256'h00000A7FF7EFEFFDFBE0000000833DFFFFADF0B9A3FFCA001BFF200F7E7AF000;
defparam sdpb_inst_5.INIT_RAM_13 = 256'h00000003BFDBFF97FFFE00000024FFFFFFEAB7CDE0BFFE4300FFF006CB02A780;
defparam sdpb_inst_5.INIT_RAM_14 = 256'hE00188017EFFDFF7FFFFE000000007FFFFFFF0E7FCB9FF808003FD842E3FEF2C;
defparam sdpb_inst_5.INIT_RAM_15 = 256'h16001F00003F6DFEFFFFDE00000078EBFFFFFA1DEFDF07FE038007F000EC7F09;
defparam sdpb_inst_5.INIT_RAM_16 = 256'hC1F803048C17BFFE3C9FF7E00000087F3FFFFFF923F6759BCC3F807F80074B75;
defparam sdpb_inst_5.INIT_RAM_17 = 256'hA213800000DFBFFFF77DFFFE10000009BFFFFFFF33BFCFF502387E07FE0179F4;
defparam sdpb_inst_5.INIT_RAM_18 = 256'h0C009E00000007FBC7A38FF7E000000B9FFFFFFFED648FFF110410F8FF740FB6;
defparam sdpb_inst_5.INIT_RAM_19 = 256'hEE6B1EF000001C53EF66E557FE0000002EFFEFFFFD2A2CDFF210B5838FFEFFF9;
defparam sdpb_inst_5.INIT_RAM_1A = 256'hEF13C83540000141FF7DE375FBE000000177FFFFFFC56068FE600457383FFFFF;
defparam sdpb_inst_5.INIT_RAM_1B = 256'h25F977884C000000FBFDEC3AAFEE00000377F7FFFFF0F7078FD6428F7987FFE5;
defparam sdpb_inst_5.INIT_RAM_1C = 256'h06E44A323E6000021FF7FFE776FF60010020F49BFFFE4EA460FF4E3F61981F79;
defparam sdpb_inst_5.INIT_RAM_1D = 256'hF4A60A58FFEB800000FFFBFF18FBFE2000006DF19CFFE0464A5620DBCCDB40C7;
defparam sdpb_inst_5.INIT_RAM_1E = 256'hA7353942DDADBC000023BBFFF37DFDE000084045017FDF000137680E81E4B018;
defparam sdpb_inst_5.INIT_RAM_1F = 256'h0F4AA03FD33775F0200279FFF80B16FE00008820000C7FE0C1807F0054C09300;
defparam sdpb_inst_5.INIT_RAM_20 = 256'h01A269C11F07DF57A0100FF7BBC4B9FFE00088002139B9E81D9827F4143D8D78;
defparam sdpb_inst_5.INIT_RAM_21 = 256'hF011E5FEDBBCD79CCE6801EFFFBD2D36FE000000080F836B419C811D829F60E7;
defparam sdpb_inst_5.INIT_RAM_22 = 256'h9F0B8BF00D196FF9661C800FCFFFFAA7FFE0000200309B0C361A202CE856659A;
defparam sdpb_inst_5.INIT_RAM_23 = 256'hEA706AEC1E15BBEE819333D4FFEFBE7B6FBE000405201FD522E3E611F9C7EB19;
defparam sdpb_inst_5.INIT_RAM_24 = 256'hBDA70F2887FCB9BFE83C3D1D3FFFFFEFC17FE000000034808100387F59C4674B;
defparam sdpb_inst_5.INIT_RAM_25 = 256'hFB6A39DA18FFE451E337E3007D6FF7ACA413FE000040070660E0038B79C53183;
defparam sdpb_inst_5.INIT_RAM_26 = 256'hAF8CB7FCD98BFFAAA17CDCEFA7FFF5FFBDA5FFC20000005C2D424C7153201404;
defparam sdpb_inst_5.INIT_RAM_27 = 256'h0CF2127FD8C8FFF81B83A50E07EFFAF7D64C7DFF00040002CD0A709EC0D180C0;
defparam sdpb_inst_5.INIT_RAM_28 = 256'h427F8263FDC58FFF95589905001CBFFDFFEF7F7FFC000000134D8F2B98B8830C;
defparam sdpb_inst_5.INIT_RAM_29 = 256'hC28B96647FFCE47FFA7C8594C00077FF7FE4ECCFFF000000000501FEB125F850;
defparam sdpb_inst_5.INIT_RAM_2A = 256'hFA48024EC7FEF627FF22F84898000F2FFFDC81939FF900000000287E462641C7;
defparam sdpb_inst_5.INIT_RAM_2B = 256'hFA30F5DD98787D5E7FE66D84D38000367FBFFD771FFF8400000003077286E61A;
defparam sdpb_inst_5.INIT_RAM_2C = 256'hEB204A67318FE372B1F8DB924F78003193FFF3CC44B3FC8000000023A14FCE3B;
defparam sdpb_inst_5.INIT_RAM_2D = 256'h000202084631FC38A08B64B4049AC0221B3FFBABE012BFC1000000019A2751C3;
defparam sdpb_inst_5.INIT_RAM_2E = 256'h80FFFE2CB8C73F40DB1C1CE3AC7186000399FFFFF43C6FFE2000004447BA32E0;
defparam sdpb_inst_5.INIT_RAM_2F = 256'h063E07714A3CE3F40CED89A5D4E3B030003B8FF7BEC851FFC8000001BFDAB603;
defparam sdpb_inst_5.INIT_RAM_30 = 256'hCBB3803B67CE38780066DBC07A9E2791801F18FFDFB0E8AFFE4000003FFFD6B0;
defparam sdpb_inst_5.INIT_RAM_31 = 256'h05CA6068E3230F0F9003AA516C67F1A82607EC4FFFEE82D77F9000002FFE5DAC;
defparam sdpb_inst_5.INIT_RAM_32 = 256'h45F1A65FD9360FC0F0001432758DFF92F71FF8B4FFF9EEB85FDF0008803FA1C5;
defparam sdpb_inst_5.INIT_RAM_33 = 256'h38F93AC7FFF99FB83F0200423EB23FFD7F9200714FF7FDE003DFC8002017F07D;
defparam sdpb_inst_5.INIT_RAM_34 = 256'hD479C7A8FC403D000FE000036C059FFFCB75AF2A1C7FF313007FFF0000097E05;
defparam sdpb_inst_5.INIT_RAM_35 = 256'h0D10988B1C005FE503FE00000CF3A3FFFECA3459064BFFF2D40BFFE080007FE0;
defparam sdpb_inst_5.INIT_RAM_36 = 256'hF1D9459E53803FFFEFFF9000000F84FFF7F46242CA3C7FF766F037FD000103FF;
defparam sdpb_inst_5.INIT_RAM_37 = 256'h7F0CA30D1A607FFFFFFFFC000128011FFDFF144CB5076BFDFDC6BBFEF000027F;
defparam sdpb_inst_5.INIT_RAM_38 = 256'h1BF4EA11036C36FFFFFFDA8000101803FFFFF9C3E1C3BA7FFF6E0FC7FE800B0E;
defparam sdpb_inst_5.INIT_RAM_39 = 256'h1FFFC72EF5E5817FFFFFFE0900012AAFFFFEFFE6548A9FD7FFE6B6C9FFA80002;
defparam sdpb_inst_5.INIT_RAM_3A = 256'h0326FE1BFE29181FFCF7DD800000047FFFD0FD7F19ABE2AFFF7F4EA01FFE0000;
defparam sdpb_inst_5.INIT_RAM_3B = 256'h0325FBF164FE6620F9D99D7104000123A0F6E3FBF87B9CFBF1E8FDBB86BFF000;
defparam sdpb_inst_5.INIT_RAM_3C = 256'h0013DFFF439830D7C71ACB8440000010800CA31FFFC47B14F1DD4FCB386FFF20;
defparam sdpb_inst_5.INIT_RAM_3D = 256'h080433FFFF060E720670013800000001000013D3FFFF6062FC3CEFEFFF0BEFF0;
defparam sdpb_inst_5.INIT_RAM_3E = 256'hB104219FFFFC1FFD95871016900000000000DDC67FFFFFE111A8E7FFBF7227FE;
defparam sdpb_inst_5.INIT_RAM_3F = 256'hFFB823B6FFFFFC1DC590FA09D7900000000D96E00FFFFFFFC78F9B3B7B673BFF;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b1;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'hFFFC005FDFDFFFF05063C780364B0000019B4CC033FFFFFFFFBD1775F7FFE377;
defparam sdpb_inst_6.INIT_RAM_01 = 256'h2FFF83012ED9B5FF0307D07E0E06CC0005EF3F800FFFFFFFFFFD3FEE7FFFDC67;
defparam sdpb_inst_6.INIT_RAM_02 = 256'hD9FFBF88EFEFBAFEFE6B5BE78080E24007BEC000047FFF81FFFFE1D71C7FFFFD;
defparam sdpb_inst_6.INIT_RAM_03 = 256'hDBBFFECC92DA0925FFC611E2F9893F8671D4F8000000180ABFFFFF1EFD53FFEF;
defparam sdpb_inst_6.INIT_RAM_04 = 256'hFBD7FFFF051096DBEFFE5F9AEF8584F8F26D580003ADD7EF40FFFFFCB7FB9FFF;
defparam sdpb_inst_6.INIT_RAM_05 = 256'hFEF77FFE7178101836FFC46AC5FC701FCBF66F200D2C92E3323BFFFFECF2A6FF;
defparam sdpb_inst_6.INIT_RAM_06 = 256'h7FFFA7FFFF230642920FF8FEDB9FADE1FFFC83981CA89F0A37A4FFFFFF66CE5F;
defparam sdpb_inst_6.INIT_RAM_07 = 256'h05FFDFFFFF90540C1920DFD81343F71C1F8FC2F49FD87800F43F705FFFFA378B;
defparam sdpb_inst_6.INIT_RAM_08 = 256'hD34FFFD7FFF6001B1039A3F958AA3F44F1F3F1BE0FF078000AA5EDC59FFFF182;
defparam sdpb_inst_6.INIT_RAM_09 = 256'h70067FF3FFDF2204EE0040FFB18F47FCD60C39AEDFD93800028560BE13DFFEEF;
defparam sdpb_inst_6.INIT_RAM_0A = 256'hD614B3FFFFFDF80187000007E2BF28FEA5A904F37FF2AF00001D97E4C03B7FFE;
defparam sdpb_inst_6.INIT_RAM_0B = 256'hFEB046AFFFFFDF00BA80A20F3E7A393FFD1FAFC77FFD07D4000693FFF9AB7FFF;
defparam sdpb_inst_6.INIT_RAM_0C = 256'hFFE588EAFFF7FFF2089C0200FFCB38A3EFBAFBFD8FFE37A200006E7FFFF7677F;
defparam sdpb_inst_6.INIT_RAM_0D = 256'hFFFF82F7D7FF7FFECFACC10017F1211C7FFE7FFE51FFD5FE40001907FFFF9E9F;
defparam sdpb_inst_6.INIT_RAM_0E = 256'hAFFFFC185F3FFFFFF0714EE537FE35124FFFFEFFB13FE2BFE100011CFFFFFEC3;
defparam sdpb_inst_6.INIT_RAM_0F = 256'h81FFFF8138FDFFCFDFA09D7B502FE704087FFBFFF2A7FDDFFF80003AC3FFFFF8;
defparam sdpb_inst_6.INIT_RAM_10 = 256'hF8CBFFF8077ECDFFFFF80F5FF7BFFE519F9FFEFFFE55FF7FFF3806071C0FFFFF;
defparam sdpb_inst_6.INIT_RAM_11 = 256'hFFCE5FFD812F353FFFBFDCEFFFF7CF88DF51FFFFFFC79FF6FFFFC000248EF7FF;
defparam sdpb_inst_6.INIT_RAM_12 = 256'hBEFCFBFFDC836FA7FFFEEB6EDF97FFF30A636FFFFFFD40F89FFFFF9006681152;
defparam sdpb_inst_6.INIT_RAM_13 = 256'h02CF840FFEC45DEB7FFFDEEF73BFFFF64877A3FFFFFF047E4DFFFD7042FAC080;
defparam sdpb_inst_6.INIT_RAM_14 = 256'h00453C6D7F8C09F23D7FEDFEFFFFDFFF8CC2D63FFFFFE567CC1FFFFFFCFE2800;
defparam sdpb_inst_6.INIT_RAM_15 = 256'h00018381C17D0C3FBBF33FCF77FFFFFFF32CDF47FFFFFC74F1CBFFFFFF87FF80;
defparam sdpb_inst_6.INIT_RAM_16 = 256'h71209C3022DD01013EBB0FBDFEF7FFFAFC64D76C3FFFFFADC428BFFFFFF18F4E;
defparam sdpb_inst_6.INIT_RAM_17 = 256'hAA02942191A1F24009DE7C3DCFFFDFFFFF922282856FFFF109A5F37FFFFFE47C;
defparam sdpb_inst_6.INIT_RAM_18 = 256'hF96028188033A200002AFFEAF5FFFFFFFFE93BD8C87FFFDD31004B3FFFFFFE2B;
defparam sdpb_inst_6.INIT_RAM_19 = 256'hFBD70002303158000001A017CCDFFEFFFF79CFBCB187FFFFB5A10D21FF9FFFF8;
defparam sdpb_inst_6.INIT_RAM_1A = 256'hFF5626160010630000002BA2BE20FFFFFFF96FBEB7D03FFFCC62015E17FDFFFF;
defparam sdpb_inst_6.INIT_RAM_1B = 256'hFFFC3C00F28188F08000017AE4D25FEDBFFC3C5CB04901FFFD8CE02644BDFFFF;
defparam sdpb_inst_6.INIT_RAM_1C = 256'hFFFFFD9D438483420000000B263F28FFFFFF0E1FF865D07F9FF080052C36EFFF;
defparam sdpb_inst_6.INIT_RAM_1D = 256'hFFFFFFFD1B00019950000001522F641FFFFFF183FEF36287F97F1C80F680995F;
defparam sdpb_inst_6.INIT_RAM_1E = 256'h18AF3FFFCB4A15F41A00000007999040FFFFFD2836ED07A801FC6010095801B1;
defparam sdpb_inst_6.INIT_RAM_1F = 256'hE4010837E07D7D52F74000000AFCC1A10FFFFF880546296EC006103D01F7800F;
defparam sdpb_inst_6.INIT_RAM_20 = 256'h050000000081E26F8C2C00004047A41468FFFFF8F0E7EAE68C02E04460333006;
defparam sdpb_inst_6.INIT_RAM_21 = 256'h000000005FC609F8BB37000080A0FEA29083FFFF891AFC0AAF4008004A06BB80;
defparam sdpb_inst_6.INIT_RAM_22 = 256'h000000003F150779DB03FC0241B77FF08202FFFFF1BF6F2A1AB6001002604A30;
defparam sdpb_inst_6.INIT_RAM_23 = 256'h700000003F19980AFDF8FFF1010C7EFBF0A047FFFE32B3FF47BFE00000C40D57;
defparam sdpb_inst_6.INIT_RAM_24 = 256'h07800000BF86D4C0C700BFFE403FFFFBFF04147FFFC2219BC02E9E00000CC1D3;
defparam sdpb_inst_6.INIT_RAM_25 = 256'hAB78000033E1869EA13E03FFF87FFFFFFFEC01A6FFFC700AE998C078000078F8;
defparam sdpb_inst_6.INIT_RAM_26 = 256'hF2E7C00001FC67D19A24F00FFF8FFFFFFFFF400D3FFF1069B6833DEF00001CAF;
defparam sdpb_inst_6.INIT_RAM_27 = 256'hFF367600007FCDD80DC84B01FFFDBFFFFFFFFF5503FFC17C94D27982780000FB;
defparam sdpb_inst_6.INIT_RAM_28 = 256'h77F427E80003F18F51E1719C01FFFFFFFFFFFF86424FF42482791F3D4F000039;
defparam sdpb_inst_6.INIT_RAM_29 = 256'h7BBC727600223E35C155FBA7700FFFFFFFFFFFFEF8C0583423881385B0E00006;
defparam sdpb_inst_6.INIT_RAM_2A = 256'h0F5FF487F610AF86B2A4EBB8B4803FF77FFFFFEFFC021C034A50607AC28E0000;
defparam sdpb_inst_6.INIT_RAM_2B = 256'h41C5FE427F871FF8D4E5C831F704007FFFFFFFFFFFFFE101ED2F978B9153F400;
defparam sdpb_inst_6.INIT_RAM_2C = 256'h033B3F8E67F136FF1A9D85C786C03004FFFFFFFFFFFFF8042F80857BF6231E00;
defparam sdpb_inst_6.INIT_RAM_2D = 256'h8693AEF49E7FBBFDD36DDB809B9D3AC01FFFFFDFFFDFBEA42CF0F84E30A4E3EE;
defparam sdpb_inst_6.INIT_RAM_2E = 256'hEF177A650EE7FEF7F02583F817FF7F290007FFDFFDFEFDD8018F2FAC382AE67F;
defparam sdpb_inst_6.INIT_RAM_2F = 256'hBFFFFF2700C23FFFFF86A45160097F326800177FF67BBFDE0433999C598CFC47;
defparam sdpb_inst_6.INIT_RAM_30 = 256'hCFFFFDE5F11260FFFFF0EB9C1C310A57546003EF84C16B09C1362EB802E8587C;
defparam sdpb_inst_6.INIT_RAM_31 = 256'hA8FFFFFC5303740FFFFC1CD8051E108C5C2D0008020800851606EFB283150203;
defparam sdpb_inst_6.INIT_RAM_32 = 256'hEA87FFFFC5F07540FFFFA1975CEB0100B702BC84000000040000BCCCB0037412;
defparam sdpb_inst_6.INIT_RAM_33 = 256'h77087FFFFC6306D40FFFF8195CF69020173A10DA6404800080000B93C3705503;
defparam sdpb_inst_6.INIT_RAM_34 = 256'h03AEC7FFFC0A3961E07FFE43907EA5B8712B71BFE7802000000009B93D000A80;
defparam sdpb_inst_6.INIT_RAM_35 = 256'h0073B847FF01837CCC03EFE0390724A4080207C4DB70001000000A1FDE800018;
defparam sdpb_inst_6.INIT_RAM_36 = 256'h100C5900A8D01CB7CAF0DEF8039278604B45110FA42FFE8260004101B9AC8000;
defparam sdpb_inst_6.INIT_RAM_37 = 256'h0066D7500428033BFE7E017700395FF345322BE90B8F2FEA000000D08F95C000;
defparam sdpb_inst_6.INIT_RAM_38 = 256'hF82DD6EB04000012BF33E04A2003CF8F4B283795CCEB37BFC03A000CD7F11413;
defparam sdpb_inst_6.INIT_RAM_39 = 256'hABF6F8F3A008000609FC5C0010003CA2339A674B5F85FCEDFED0E00281F78881;
defparam sdpb_inst_6.INIT_RAM_3A = 256'hCBB3B09BD7000001EF9E4DE0000003E84FE5E42FA2FC89F02FEDE5BA7EFFF8AE;
defparam sdpb_inst_6.INIT_RAM_3B = 256'h488B752FD84000007CB80E4D0000007E5641A97E7C868D3E7EEFFFFF7FFFFECD;
defparam sdpb_inst_6.INIT_RAM_3C = 256'h837D9DAF0E28000007A208E1E0000001C6BFDD46EF40BCE2EA0A7FFB4BFE7F78;
defparam sdpb_inst_6.INIT_RAM_3D = 256'hE809F978552780010FE464329C000020FF34236233CB21B60FC8E03FFFFFF7FF;
defparam sdpb_inst_6.INIT_RAM_3E = 256'hDF40C50534B718000BFEB7FE19EC0A404FF1AF9A6FCE5CD1E9ECF685FFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3F = 256'hFFF007150698A70931DFC307DD9FF88093FF8CBB05F6934318FE1C107FFFDFFF;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b1;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'h200CA7CFBFFFFFFFFF20100000001BFFFFFFFFFFFF7FFDFDFFFFFFFFFFFFFE84;
defparam sdpb_inst_7.INIT_RAM_01 = 256'hE000EEBFFDFFFFFFFFE2000C000009AFFFFFFFFFFFFF6FE3AFFFFFFFFFFFFFF8;
defparam sdpb_inst_7.INIT_RAM_02 = 256'hFF0077BFFFFFFFFFFFFD0002E0000002BF7FFFFF7B860C03C5DFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_03 = 256'hFFF880FFFFFFFFFFFFFA0800FFC00000637EFFFA82028004861CFB7FFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_04 = 256'hFFFFC1F9FFFFFFFFFFFF84003FFE00004010F05C9000000011C4407FFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_05 = 256'hFFFFF90DFFFFFFFFFFFFFE0001FFE1000100772B00B200000115401FFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_06 = 256'hFFFFFFE1FFEFFFFFFFFFEF00001BFE700000473A1864000000003806EFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_07 = 256'hFFFFFFFF7FFFFFFFFFFFFFF8206FCF0FD0040DBF9A0600000000906E5A7FFFFF;
defparam sdpb_inst_7.INIT_RAM_08 = 256'hFFFFFFFFF7FFFFFFFFFFFFFE8003FD5FFF001C17FA50000000000100777FFFFF;
defparam sdpb_inst_7.INIT_RAM_09 = 256'hFFFFFFFFFEFFEDFFFFFFFFFFFC02FFF7FFFFFEE9FF7B06004000800800BDFFFF;
defparam sdpb_inst_7.INIT_RAM_0A = 256'hFFFFFFFFFFFFEFFFBFFFFFFFFE401FFDDBFFB7FFB77FB480540B0000417BF6FB;
defparam sdpb_inst_7.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE822FFEAEFEFDFFFFFFF8000002350002FEDAF;
defparam sdpb_inst_7.INIT_RAM_0C = 256'h71FEFF9FFFFFF7FFFFFFFFFFFFFF23C9F8FF97FF3FFFFDF0000000B500006EED;
defparam sdpb_inst_7.INIT_RAM_0D = 256'hEFFFFFFFFFFFFFFFFFF7FFFFFFFF5C7EAB3FFF3FFCFFFFFE00007C100081046F;
defparam sdpb_inst_7.INIT_RAM_0E = 256'h6FDFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFA8FFFDBFF5FFFFFE0103A3C28E8004F;
defparam sdpb_inst_7.INIT_RAM_0F = 256'hA7DBFF3FFFFFFFFFF7FFFFFFFFFFFFADFFCAFFF9B7FDFFFFFA000D0C7000B023;
defparam sdpb_inst_7.INIT_RAM_10 = 256'h00CE1EF29FFFFBFFFFFFFFFFFFFFFFFFBFF8EBFDBEFB3FFFFF000387F7000100;
defparam sdpb_inst_7.INIT_RAM_11 = 256'h00077FFFFBFFFDFFFFFFFFFFFFFFFFFFF8FFBEA7D7F2DEFFFFF4402185CA0000;
defparam sdpb_inst_7.INIT_RAM_12 = 256'h00000A7FF7EFEFFDFBFFFFFFFFFFFFFFFFA7E7FAC9FFCFEFFFFF200D8F8DF000;
defparam sdpb_inst_7.INIT_RAM_13 = 256'h00000003BFDBFF97FFFFFFFFFFFFFFFFFFEF817FE17FFEFFFFFFF006FC3D5B80;
defparam sdpb_inst_7.INIT_RAM_14 = 256'hE00188017EFFDFF7FFFFFFFFFFFFFFFFFFFFF89FFC79FF5FEFFFFD842F8A105C;
defparam sdpb_inst_7.INIT_RAM_15 = 256'hEE001F00003F6DFEFFFFDFFFFFFFFFFFFFFFFFEBFFE037F17E7FFFF000F4007A;
defparam sdpb_inst_7.INIT_RAM_16 = 256'h2EB803048C17BFFE3C9FF7FFFFFFFFFFFFFFFFFFBBF071D83FE07FFF8007BC9D;
defparam sdpb_inst_7.INIT_RAM_17 = 256'hC8EB800000DFBFFFF77DFFFFFFFFFFFFFFFFFFFDF6DE2FF7ED3A01FFFE017C48;
defparam sdpb_inst_7.INIT_RAM_18 = 256'hC777EE00000007FBC7A38FF7FFFFFFFFFFFFFFFFFF5D33FF5AFC3007FF740FDE;
defparam sdpb_inst_7.INIT_RAM_19 = 256'hF53DCBF000001C53EF66E557FFFFFFFFFFFFFFFFFFBDE3DFF5EFAF807FFEFFFE;
defparam sdpb_inst_7.INIT_RAM_1A = 256'hFFD77F9F40000141FF7DE375FBFFFFFFFFFFFFFFFFF39F98FE2BFFFF07FFFFFF;
defparam sdpb_inst_7.INIT_RAM_1B = 256'hA13E224FBC000000FBFDEC3AAFEFFFFFFFFFFFFFFFFFEBFFCFC1BF3FF87FFFFA;
defparam sdpb_inst_7.INIT_RAM_1C = 256'hCE5070998EE000021FF7FFE776FF7FFFFFFFFFFFFFFFFFFBEBBC3FFFFF87FFF1;
defparam sdpb_inst_7.INIT_RAM_1D = 256'h6E1F6F84EFA7800000FFFBFF18FBFFDFFFFFFFFFFFFFFFFFFEAB8FF97E38BFFA;
defparam sdpb_inst_7.INIT_RAM_1E = 256'hC8B29CEC07EF9C000023BBFFF37DFDFFFFFFFFFFFFFFFFFFDFF89FFF77E38FFF;
defparam sdpb_inst_7.INIT_RAM_1F = 256'hF38CFAECA4BF3CF0200279FFF80B16FFFFFFFFFFFFFFFFFF1F7E80FF3F8CB0FF;
defparam sdpb_inst_7.INIT_RAM_20 = 256'hFE0339EAFCBDED77A0100FF7BBC4B9FFFFFFFFFFFFDFF3FFE267C00FF7FA8B07;
defparam sdpb_inst_7.INIT_RAM_21 = 256'h0FE7A0008FB1C7FFFE6801EFFFBD2D36FFFFFFFFFFF77FBFFE26FFA2BE1F30A0;
defparam sdpb_inst_7.INIT_RAM_22 = 256'h80F4BF4FF1318F7FFDFC800FCFFFFAA7FFFFFFFFFFFFA381FBE387F50FA3E980;
defparam sdpb_inst_7.INIT_RAM_23 = 256'hC60F82EBFFE1B06AFA70B3D4FFEFBE7B6FBFFFFFFFFFE07D1D1C389FD7BD9D5B;
defparam sdpb_inst_7.INIT_RAM_24 = 256'hD560F10D7FFF09E31E403DFD3FFFFFEFC17FFFFFFFFFFF07F3FBC08DFB31FDBD;
defparam sdpb_inst_7.INIT_RAM_25 = 256'hFE660618D7FFF9DE10E87CFDFD6FF7ACA413FFFFFFFFFB9D5F3E7C0CAB7CFFCF;
defparam sdpb_inst_7.INIT_RAM_26 = 256'hDFCC7001657FFFC48EC30FB015FFF5FFBDA5FFFDFFFFFFA0D5E28B81E597EBFF;
defparam sdpb_inst_7.INIT_RAM_27 = 256'hE6FC0E001D07FFFE9B760391F86FFAF7D64C7DFEFFFBFFF9089960E0F72E1FFF;
defparam sdpb_inst_7.INIT_RAM_28 = 256'hBFEF81E001657FFFEA873B7AFFE2FFFDFFEF7F7FE3FFFFFFEA68AF2C1EC77DF7;
defparam sdpb_inst_7.INIT_RAM_29 = 256'h789DBE1C001413FFFCA5787F3FFF97FF7FE4ECCFFEFFFFFFFFF881FE41C617FF;
defparam sdpb_inst_7.INIT_RAM_2A = 256'hFD3BCFC1C000E09FFFD4979CE7FFF0DFFFDC81939FE6FFFFFFFFC07FE0387F7F;
defparam sdpb_inst_7.INIT_RAM_2B = 256'hE5F67C7C780789D5FFFA1379FF7FFFCFFFBFFD771FFE7BFFFFFFFE07AE0707FB;
defparam sdpb_inst_7.INIT_RAM_2C = 256'hEB3FDFE70F801C784FFF5AAF9E87FFCEEFFFF3CC44B3E37FFFFFFFDDDC47F03F;
defparam sdpb_inst_7.INIT_RAM_2D = 256'h00017FF841F003C3827F8F89F9E13FDDE7FFFBABE012BE3EFFFFFFFE5FF03E03;
defparam sdpb_inst_7.INIT_RAM_2E = 256'h800005FEB83F00BF0FD3E7141F94B9FFFC77FFFFF43C6FE1DFFFFFBBBB840100;
defparam sdpb_inst_7.INIT_RAM_2F = 256'h7E01F86FDE03E00BF1CA81D9A3FD09CFFFC57FF7BEC851FE37FFFFFE406CB783;
defparam sdpb_inst_7.INIT_RAM_30 = 256'h20707FC379C1F807FF89BC033C7FCD1E7FE0B7FFDFB0E8AFE1BFFFFFC002CB38;
defparam sdpb_inst_7.INIT_RAM_31 = 256'h02461FFF00C0FF006FFC9C33575FFE90D9F81B3FFFEE82D77E6FFFFFD0002DCF;
defparam sdpb_inst_7.INIT_RAM_32 = 256'h802F61FFFEEBFFC00FFFE4F060E3FFE620E00693FFF9EEB85FE0FFF77FC002D6;
defparam sdpb_inst_7.INIT_RAM_33 = 256'h8C07963FFFF81FB800FDFF95F769FFFE59C1FFC33FF7FDE003DE37FFDFE80076;
defparam sdpb_inst_7.INIT_RAM_34 = 256'hF8802D67FC400000001FFFFC5CB07FFFF2C583C8F3FFF313007FE0FFFFF68007;
defparam sdpb_inst_7.INIT_RAM_35 = 256'h0E277B26FC0000000001FFFFF0FCDFFFFF17ADD12B3FFFF2D40BFE1F7FFF8000;
defparam sdpb_inst_7.INIT_RAM_36 = 256'h01E33852CF80000000006FFFFFF003FFF7F8A4E2C1FBFFF766F037E2FFFEFC00;
defparam sdpb_inst_7.INIT_RAM_37 = 256'h800F30A349E00000000003FFFFFFFEFFFDFFE6FB56FE1FFDFDC6BBFF0FFFFD80;
defparam sdpb_inst_7.INIT_RAM_38 = 256'hE400F388891C00000000257FFFFFFFFFFFFFFE1ABFDFDDFFFF6E0FC7E17FF4F1;
defparam sdpb_inst_7.INIT_RAM_39 = 256'hE00007CBCB238000000001F6FFFFFFFFFFFEFFF866A7EBEFFFE6B6C9FE57FFFD;
defparam sdpb_inst_7.INIT_RAM_3A = 256'hFCD9001C6518F8000308227FFFFFFFFFFFFFFD7FE1CEAFB7FF7F4EA01FE1FFFF;
defparam sdpb_inst_7.INIT_RAM_3B = 256'hFCDA040178FE1E200626628EFBFFFFFFFFF8FFFBFF83CCFBC7E8FDBB86BE0FFF;
defparam sdpb_inst_7.INIT_RAM_3C = 256'hFFEC200003E00FD7C0E5347BBFFFFFFFFFFF773FFFFF82856BBD4FCB386FE0DF;
defparam sdpb_inst_7.INIT_RAM_3D = 256'hF7FBCC000007F1FDFE0FFEC7FFFFFFFFFFFF8557FFFFFF8C7F7FEFEFFF0BEE0F;
defparam sdpb_inst_7.INIT_RAM_3E = 256'h4EFBDE6000001FFEC860EFE96FFFFFFFFFFF3C41FFFFFFFE656BFFFFBF7227E1;
defparam sdpb_inst_7.INIT_RAM_3F = 256'hE047DC490000001DE6AA05F6106FFFFFFFF14A9FFFFFFFFFFB2EFF7B7B673BFE;

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[30:0],sdpb_inst_8_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_8.READ_MODE = 1'b1;
defparam sdpb_inst_8.BIT_WIDTH_0 = 1;
defparam sdpb_inst_8.BIT_WIDTH_1 = 1;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_8.RESET_MODE = "SYNC";
defparam sdpb_inst_8.INIT_RAM_00 = 256'hFE03FFA0202000005DDAE07FCDB0FFFFFE175E3FFFFFFFFFFFD976B3F7FFE377;
defparam sdpb_inst_8.INIT_RAM_01 = 256'h2FE07CFED1264A00039A9A01F1F923FFFA58007FFFFFFFFFFFFE0FFCFFFFDC67;
defparam sdpb_inst_8.INIT_RAM_02 = 256'hD9FE4077101045010075A6207F7F1D3FF8083FFFFFFFFFFFFFFFF8472EFFFFFD;
defparam sdpb_inst_8.INIT_RAM_03 = 256'hDBBFE1336D25F6DA00073D760676C0798E1A87FFFFFFFFF37FFFFFC2FBF7FFEF;
defparam sdpb_inst_8.INIT_RAM_04 = 256'hFBD7FE00FAEF692410006765607A3B07CD83C7FFFC163F0FFFBFFFFE57FFFFFF;
defparam sdpb_inst_8.INIT_RAM_05 = 256'hFEF77FE18E87EFE7C90006352C038BE0300000DFF04B32C3FC47FFFFF3FBCDFF;
defparam sdpb_inst_8.INIT_RAM_06 = 256'h7FFFA7FE00DCF9BD6DF000D31580527E01812867E17980F46AAABFFFFF9FF7EF;
defparam sdpb_inst_8.INIT_RAM_07 = 256'hFBFFDFFFE06FABF3E6DF201C0DA008E1E050220B60EE07FF7CEF3ADFFFFDFEBB;
defparam sdpb_inst_8.INIT_RAM_08 = 256'h6EDFFFD7FE09FFE4EFC65C01F1F600BB3E0A0481F04F07FFFDE9FDDF9FFFEFBC;
defparam sdpb_inst_8.INIT_RAM_09 = 256'hEF39FFF3FFE0DDFB11FFBF0036F6C00329F305A1201F87FFFD85018087DFFF7F;
defparam sdpb_inst_8.INIT_RAM_0A = 256'hFBCB07FFFFFE07FE78FFFFF80391D8015A4ED0788001A0FFFFD5FFFF543B7FFB;
defparam sdpb_inst_8.INIT_RAM_0B = 256'hFFDB887FFFFFE0FF457F5DF0C05E530002E0B4510000D02BFFF80FFFFEE97FFF;
defparam sdpb_inst_8.INIT_RAM_0C = 256'hFFFEFB17FFF7FE0DF763FDFF000F12E010450108C000845DFFFF17FFFFFA4B7F;
defparam sdpb_inst_8.INIT_RAM_0D = 256'hFFFFD4040FFF7FE130533EFFE801DCB40001800058002B01BFFFE83FFFFFF65F;
defparam sdpb_inst_8.INIT_RAM_0E = 256'h0FFFFEA0A07FFFFE0F8EB11AC80036A8C000010039000C801EFFFE03FFFFFF61;
defparam sdpb_inst_8.INIT_RAM_0F = 256'hF8FFFFF4050FFFCFE05F6284AFD006169800040000A00100007FFFC93FFFFFFD;
defparam sdpb_inst_8.INIT_RAM_10 = 256'hFECFFFFFA8423FFFFE07F0A00840007E6D8001000034000800C7F9F883FFFFFF;
defparam sdpb_inst_8.INIT_RAM_11 = 256'hFFFEBFFFFD40CAFFFFE023100008300FE2B00000000B801800003FFFCCFFFFFF;
defparam sdpb_inst_8.INIT_RAM_12 = 256'hFFFF3BFFFFE0B4DBFFFE148120680003B5A70000000170000000006FF967FFFF;
defparam sdpb_inst_8.INIT_RAM_13 = 256'hFFFFFE9FFFFF40149FFFE1108C4000087F2B600000001A006C00028FBD163FFF;
defparam sdpb_inst_8.INIT_RAM_14 = 256'hFFFFFFBAFFFFF00062FFFE01000020000E41AE00000005200A8000000300E3FF;
defparam sdpb_inst_8.INIT_RAM_15 = 256'hFFFFFFFCCFFFFFC80C27FFE08800000003CC8AC0000000340108000000780F1F;
defparam sdpb_inst_8.INIT_RAM_16 = 256'h2FFFFFFFD9FFFFFE8040BFFE01080005007AD25C0000000BC03B8000000E701D;
defparam sdpb_inst_8.INIT_RAM_17 = 256'h3EFFFFFFFF8FFFFFF44101FFE0002000001C1A19800000013807900000001B85;
defparam sdpb_inst_8.INIT_RAM_18 = 256'h02A7FFFFFFD0FFFFFFA05817FE000000000E3544B800000033005300000001D4;
defparam sdpb_inst_8.INIT_RAM_19 = 256'h04173FFFFFFC27FFFFFD94303FE001000002A5FFF780000006200AE000000007;
defparam sdpb_inst_8.INIT_RAM_1A = 256'h00A8BEFFFFFFB8FFFFFFC81E55FE00000001EFDCC1300000005E01C600000000;
defparam sdpb_inst_8.INIT_RAM_1B = 256'h0003C4CFFFFFF00FFFFFFE65820FE01240001C5E71E70000000B603AC0000000;
defparam sdpb_inst_8.INIT_RAM_1C = 256'h0000021B7FFFFC0DFFFFFFF30581FE0000000E1FCD27300000006806FC000000;
defparam sdpb_inst_8.INIT_RAM_1D = 256'h000000012A7FFE7A0FFFFFFE91400BE000000103ED92518000001980C1800000;
defparam sdpb_inst_8.INIT_RAM_1E = 256'h000000000E3FEA1481FFFFFFF980701E0000003834C70298000001500C780000;
defparam sdpb_inst_8.INIT_RAM_1F = 256'h0000000000449BBEFE3FFFFFF50C0020E000000B079EE025C0000033019B8000;
defparam sdpb_inst_8.INIT_RAM_20 = 256'h0000000000C1265BFB63FFFFBFB8200856000000C0F3EE04DC00000720387000;
defparam sdpb_inst_8.INIT_RAM_21 = 256'h000000005FE1CD9C0090FFFF7F5F0382902000000D1CFD0012C000005E075780;
defparam sdpb_inst_8.INIT_RAM_22 = 256'h000000003FE1FB7E568803FDBE4880188000000001DF9F9600AE0000076074F0;
defparam sdpb_inst_8.INIT_RAM_23 = 256'hF00000003FE07FF8FFF8000EFEF38104F07000000039F7EEC056E000008C0E2F;
defparam sdpb_inst_8.INIT_RAM_24 = 256'hDF800000BFF89AFF6F000001BFC0000407140000000347DB9C108E00000FC1EA;
defparam sdpb_inst_8.INIT_RAM_25 = 256'hD4F8000033FE15DFFC7E000007800000002C006000005372E907E5F80000C8FE;
defparam sdpb_inst_8.INIT_RAM_26 = 256'hFD5FC00001FF85703FC4F00000700000000140040000185FDAA0E0DF000017AF;
defparam sdpb_inst_8.INIT_RAM_27 = 256'hFFDDF600007FF1BCF3675B000002400000000D80C000027694CA0879F800001B;
defparam sdpb_inst_8.INIT_RAM_28 = 256'hD7F99FE80003FE14C608F9DC0000000000000037A80000AFE27F01003F00003D;
defparam sdpb_inst_8.INIT_RAM_29 = 256'h61BF89F600223FC6B4EA73CFF0000000000000008600002FBB88506C17E00007;
defparam sdpb_inst_8.INIT_RAM_2A = 256'h0E7FF9BFF610AFF8D31B1587EE80000880000010000000048C303004327E0000;
defparam sdpb_inst_8.INIT_RAM_2B = 256'h41FBFFA9FF871FFF19C3B7C938FC00000000000000000001962385802B4FF400;
defparam sdpb_inst_8.INIT_RAM_2C = 256'h033CDFF19FF136FFE336FE3C409DF00000000000000000003040F59B4168FE00;
defparam sdpb_inst_8.INIT_RAM_2D = 256'h8693DDFF09FFBBFDFC764FEF240427C000000000000000042E02F9CE70939FEE;
defparam sdpb_inst_8.INIT_RAM_2E = 256'hEF177EDFF19FFEF7FFC6BEFEE841B77D000000000000000001C02F8B4928F1FF;
defparam sdpb_inst_8.INIT_RAM_2F = 256'hFFFFFFCCFF71FFFFFFF8CE195FF284CF2800000000000000043D8A1C458C893F;
defparam sdpb_inst_8.INIT_RAM_30 = 256'h3FFFFDF8CFE31FFFFFFF0DE3BBEEF58952E00000000000000137FE0040E83A13;
defparam sdpb_inst_8.INIT_RAM_31 = 256'h47FFFFFFB0FC13FFFFFFE080FEA3FF33A29F0000000000000006FBB1038507A5;
defparam sdpb_inst_8.INIT_RAM_32 = 256'h547FFFFFF84F813FFFFFFE1B07F4FCFFFDE8BC84000000000000BF3C00057438;
defparam sdpb_inst_8.INIT_RAM_33 = 256'h11E7FFFFFFA8F813FFFFFFE1B3F77BFFEFBFEA7A6400800000000BE3C3700102;
defparam sdpb_inst_8.INIT_RAM_34 = 256'h000E3FFFFFF286871FFFFFFC1BB6B0838F3BFE9EFF802000000009BEBD000700;
defparam sdpb_inst_8.INIT_RAM_35 = 256'h000DA7FFFFFE288163FFFFFFC1BCA08897C287F9A170001000000A1FE3800008;
defparam sdpb_inst_8.INIT_RAM_36 = 256'h000224FFFFFFE2881A0FFFFFFC19A1FE223A100FC6DFFE8260004101BEBC8000;
defparam sdpb_inst_8.INIT_RAM_37 = 256'h00012D4FFFFFFC080321FFFFFFC1BB08BC01C2000D143FEA000000D08FE3C000;
defparam sdpb_inst_8.INIT_RAM_38 = 256'h00002210FFFFFFE1802E1FFFFFFC0A5020FD184A00D71CFFC03A000CD7FE4C00;
defparam sdpb_inst_8.INIT_RAM_39 = 256'h800007E49FFFFFF8580743FFFFFFC0D1038DE620A006040DFED0E00281F7F260;
defparam sdpb_inst_8.INIT_RAM_3A = 256'h56E80EF450FFFFFE0680641FFFFFFC0ECE7CF0A8DD00D8219FFDE5BA7EFFFF39;
defparam sdpb_inst_8.INIT_RAM_3B = 256'h8D3A55CFAA3FFFFF816809C2FFFFFF806247207E03790A2F4B7FFFFF7FFFFFF1;
defparam sdpb_inst_8.INIT_RAM_3C = 256'hFC6A7BA31267FFFFF83080A81FFFFFFE0711ED26EABF4081F30DFFFB4BFE7FFF;
defparam sdpb_inst_8.INIT_RAM_3D = 256'hFFF122DB4E4C7FFEF0062C3683FFFFDF00397D0FB31EDE383F68FFFFFFFFF7FF;
defparam sdpb_inst_8.INIT_RAM_3E = 256'hFFFF0646350507FFF400F77FC813F5BFB001CA1DD7B2132127F0F6FFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3F = 256'hFFFFF819AC5260F6CE200F4FF680077F6C000F28BF601FBC047F4C0FFFFFFFFF;

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[29:0],sdpb_inst_9_dout[3:2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[15],ada[14],ada[13]}),
    .BLKSELB({adb[15],adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_9.READ_MODE = 1'b1;
defparam sdpb_inst_9.BIT_WIDTH_0 = 2;
defparam sdpb_inst_9.BIT_WIDTH_1 = 2;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_9.RESET_MODE = "SYNC";
defparam sdpb_inst_9.INIT_RAM_00 = 256'h5595556555403E904B11CFF4BF1A97B26032ECAFE9C0F00F0AABFFFFFFFFFFFB;
defparam sdpb_inst_9.INIT_RAM_01 = 256'hBBEEAAFBAAAA95503E53A96B1BC1559AA99595555540D8647F9BE5F055556559;
defparam sdpb_inst_9.INIT_RAM_02 = 256'h5555595555555003E93471D7FF8C6A003FF3E461BFE785F00D26AAFEBFABBFEF;
defparam sdpb_inst_9.INIT_RAM_03 = 256'hEEBAAAABABBEAAA95503EEA6AAFC0555A999595555550FF479BE4335C0555559;
defparam sdpb_inst_9.INIT_RAM_04 = 256'h556655555555555500FE9376FDBFFA4B7C35B616BDFFA301F00C6E5AABEFAAFB;
defparam sdpb_inst_9.INIT_RAM_05 = 256'hEBABEEAEAEAAEAEAAA555400CF3001559555965555555403BD91BE7F19C15555;
defparam sdpb_inst_9.INIT_RAM_06 = 256'h565555555555555555000FA53B1BE701ACFF0F4C9FAD6F91C3C0DDC59ABAABEA;
defparam sdpb_inst_9.INIT_RAM_07 = 256'hEAAAAEAAAEAAAAAAAAAA99544500000555565556555555554F9336FE7BFEC155;
defparam sdpb_inst_9.INIT_RAM_08 = 256'h15555555555555555554000FFA5371AB843CBCF034D66D1A4CC2C40C6916AAAA;
defparam sdpb_inst_9.INIT_RAM_09 = 256'hAAAAAAAAAAAAAAAAAA9AAAA55555055455555555555555554403E01BFE6306C5;
defparam sdpb_inst_9.INIT_RAM_0A = 256'hC1145555555555555555550003FFE97A6BB153E53C33F060565B0014438E0AAA;
defparam sdpb_inst_9.INIT_RAM_0B = 256'hAAAA9AAABAAAAAAAAAA6A9A5595555554555565595555555554400FEBCFE0B67;
defparam sdpb_inst_9.INIT_RAM_0C = 256'hBB05545555555555555555151103CFFEA49B81553B250E8861AA58181500E1CA;
defparam sdpb_inst_9.INIT_RAM_0D = 256'h05AAAAAAA9AAAA6AA5AAA5A66A6A59655555555555555145555500003FCC0E38;
defparam sdpb_inst_9.INIT_RAM_0E = 256'h59EC01055554155555105515045040003FF94DCE1942F0F1232B597735514039;
defparam sdpb_inst_9.INIT_RAM_0F = 256'h3BC55AAAAAAAA9AAAAAAAAA6595695665555555555555515401154000000000E;
defparam sdpb_inst_9.INIT_RAM_10 = 256'h03A1B000050505541510114554555500000CFFA4E3AE543D80CACAD571055540;
defparam sdpb_inst_9.INIT_RAM_11 = 256'h403F856AAAAAAA6AA95A95996595655555555555555554114000101000000000;
defparam sdpb_inst_9.INIT_RAM_12 = 256'h0003FFF000000014154004154105105400011000FE92259543D68AFA853C9515;
defparam sdpb_inst_9.INIT_RAM_13 = 256'h450034055669AAAAAA6955665555565555595555555555555000000000440000;
defparam sdpb_inst_9.INIT_RAM_14 = 256'h0000000000000040000000000000000400410100003FA4EE7854E4EBE1EF9655;
defparam sdpb_inst_9.INIT_RAM_15 = 256'h155510ECC1555AA9A96999555555555555555555555515514000003000000400;
defparam sdpb_inst_9.INIT_RAM_16 = 256'h000C0000000000000000000000010000D4400045054000FE9D97A50FC5CC384F;
defparam sdpb_inst_9.INIT_RAM_17 = 256'hA0754501ABC555A5595555665555555555555555555515555400000000000000;
defparam sdpb_inst_9.INIT_RAM_18 = 256'h000000000000300000000CC00003000000000000545414000FA4996850520602;
defparam sdpb_inst_9.INIT_RAM_19 = 256'h8A0551054192C15559565655955555555555515555551454554100000C000000;
defparam sdpb_inst_9.INIT_RAM_1A = 256'hC3000C0F0C3F0000030303000000003000000000000055514100FA4871D4F12A;
defparam sdpb_inst_9.INIT_RAM_1B = 256'h54FA44034040AF055555559555555555555550005500501550444000300FCF03;
defparam sdpb_inst_9.INIT_RAM_1C = 256'hCFCFCCFFFFFFF000F0CCF0F00000F03F300000000C0005455551440FA780544E;
defparam sdpb_inst_9.INIT_RAM_1D = 256'h23F50A5453003F2B01555555556555554055500440040040001000000003CCC3;
defparam sdpb_inst_9.INIT_RAM_1E = 256'hF3FFFFFFFFFFFFFC0FF0CCFCCFC0FC0FFCC3333C000000011155555000E9370B;
defparam sdpb_inst_9.INIT_RAM_1F = 256'h215A7D99515040016B04555555545555001010000000000000004000003F0FFF;
defparam sdpb_inst_9.INIT_RAM_20 = 256'hFFCFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFCFF330000054555555103E92;
defparam sdpb_inst_9.INIT_RAM_21 = 256'hE5E1105B5E044C7C386805555555555545000000000000000000000000003FFF;
defparam sdpb_inst_9.INIT_RAM_22 = 256'hFFFBFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF30000111555555403;
defparam sdpb_inst_9.INIT_RAM_23 = 256'h403E4E22E5BF201BFBE37C0155555055545100000000000000000000000003FF;
defparam sdpb_inst_9.INIT_RAM_24 = 256'hFFFAFFFBFBFBFBFFFFFFFFFBFFFFFFFFFFFFFBFFEBFFFFCFCFCC000115555555;
defparam sdpb_inst_9.INIT_RAM_25 = 256'h555403E5E35F3E8BFEA7A2B005554555055050000C00000C0CC30300300C03FF;
defparam sdpb_inst_9.INIT_RAM_26 = 256'hFFFFBFEEFEBBEAAAFAFEBFFFFFFEFFFFBEFBFBEBFBBAFFFFFFFFF00000155555;
defparam sdpb_inst_9.INIT_RAM_27 = 256'h55555500FA4E715F04A0471AFC00515144004511433FF0C0FFCFFC3C0F3F000F;
defparam sdpb_inst_9.INIT_RAM_28 = 256'h3FFFFAAAAAAAAABABAAEAFAEFEFABEBABAAFEAAAEAAEAEBEBEAFFFFC00001455;
defparam sdpb_inst_9.INIT_RAM_29 = 256'h55555555500FE42218BBB2EB06C04505500000110003FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2A = 256'hFFFFBBAEBAAAAAAAB9AAAAAABAABAAAAAAAAAAAAAAAAEAAAAAAFAAFFFFC00001;
defparam sdpb_inst_9.INIT_RAM_2B = 256'h00055595555400FE53789C0660DB01055150100000000CFBFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2C = 256'hFFFBBFEAAA9AAAAAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABFFFFC0;
defparam sdpb_inst_9.INIT_RAM_2D = 256'hF00001555555551003E94E83BCB06FC015400400040000CFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_9.INIT_RAM_2E = 256'hFFFBBAEEAAAAA9566AAAA66AAAAAAAAAAAAAAAAA9AAAAA569AA566AAAAABBFFF;
defparam sdpb_inst_9.INIT_RAM_2F = 256'hFFF0C0005455555555503FA943F05AFC011404400000000333FFEEFFFBFEFEEA;
defparam sdpb_inst_9.INIT_RAM_30 = 256'hEAAAAFEAAA9965995655695A655AA999AA6AAAAA5956A65965555669566AAAAB;
defparam sdpb_inst_9.INIT_RAM_31 = 256'hA6EBFFF00001555555555503FBAAAAABF0041440000000000FFEFEEBBFAABABF;
defparam sdpb_inst_9.INIT_RAM_32 = 256'hAAAAAAAAAA95655555555559555555559A5595555655555555555555565559AA;
defparam sdpb_inst_9.INIT_RAM_33 = 256'h00000000000000000000000000000000000000000000000000000002AAAFAAAA;

SDPB sdpb_inst_10 (
    .DO({sdpb_inst_10_dout_w[30:0],sdpb_inst_10_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_10.READ_MODE = 1'b1;
defparam sdpb_inst_10.BIT_WIDTH_0 = 1;
defparam sdpb_inst_10.BIT_WIDTH_1 = 1;
defparam sdpb_inst_10.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_10.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_10.RESET_MODE = "SYNC";
defparam sdpb_inst_10.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFF20100000001BFFFFFFFFFFFF7FFDFDFFFFFFFFFFFFFFF8;
defparam sdpb_inst_10.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFE20008000009AFFFFFFFFFFFFF6FE3AFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFD0003E0000002BF7FFFFF7B860C03C5DFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFA0800FFC00000637EFFFA82028004861CFB7FFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFF84003FFF00004010F05C9000000011C4407FFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFE0003FFFF000100772B00B200000115401FFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFEF0000FBFBF80000473A1864000000003806EFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFF8206EEECFF0040DBF9A0600000000906E5A7FFFFF;
defparam sdpb_inst_10.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE8007FBD3FF801C17FA50000000000100777FFFFF;
defparam sdpb_inst_10.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC03FFECFFF7FEE9FF7B06004000800800BDFFFF;
defparam sdpb_inst_10.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE401FFDFBFEB7FFB77FB480540B0000417BF6FB;
defparam sdpb_inst_10.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE826FFB26FBFDFFFFFFF8000002350002FEDAF;
defparam sdpb_inst_10.INIT_RAM_0C = 256'h71FEFF9FFFFFFFFFFFFFFFFFFFFF23D9ECF994FF7FFFFDF0000000B500006EED;
defparam sdpb_inst_10.INIT_RAM_0D = 256'hEFFFFFFFFFFFFFFFFFFFFFFFFFFF5C3F6BBFE7BFFFFFFFFE00007C100081046F;
defparam sdpb_inst_10.INIT_RAM_0E = 256'h6FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDE7FFCFFF7FFFFFE01039EC28E8004F;
defparam sdpb_inst_10.INIT_RAM_0F = 256'hA7DBFF3FFFFFFFFFFFFFFFFFFFFFFFAFFFD0FFED67EBFFFFFA000D9A7000B023;
defparam sdpb_inst_10.INIT_RAM_10 = 256'h00CE1EF29FFFFBFFFFFFFFFFFFFFFFFFBFFF7BFD7DBB7FFFFF0003F4A7000100;
defparam sdpb_inst_10.INIT_RAM_11 = 256'h00077FFFFBFFFDFFFFFFFFFFFFFFFFFFF7FF5F6767FE6EFFFFF4403D540A0000;
defparam sdpb_inst_10.INIT_RAM_12 = 256'h00000A7FF7EFEFFDFBFFFFFFFFFFFFFFFFBBF9FDCDFFBBEFFFFF200FFC1FB000;
defparam sdpb_inst_10.INIT_RAM_13 = 256'h00000003BFDBFF97FFFFFFFFFFFFFFFFFFEFE67FFD3FFC3FFFFFF006E7CFFD80;
defparam sdpb_inst_10.INIT_RAM_14 = 256'hE00188017EFFDFF7FFFFFFFFFFFFFFFFFFFFB9CFFC59FF6BEFFFFD842F79FFDC;
defparam sdpb_inst_10.INIT_RAM_15 = 256'h9E001F00003F6DFEFFFFDFFFFFFFFFFFFFFFFFFBFFD9E7EB3EFFFFF000FB7FD9;
defparam sdpb_inst_10.INIT_RAM_16 = 256'h007803048C17BFFE3C9FF7FFFFFFFFFFFFFFFFDFDBF7769BFB9FFFFF8007DFEB;
defparam sdpb_inst_10.INIT_RAM_17 = 256'h010D800000DFBFFFF77DFFFFFFFFFFFFFFFFFFFFFA7EDFEA5FFCFFFFFE017EFC;
defparam sdpb_inst_10.INIT_RAM_18 = 256'h4C840E00000007FBC7A38FF7FFFFFFFFFFFFFFFFFF1B9BFF2BF0BFFFFF740FEF;
defparam sdpb_inst_10.INIT_RAM_19 = 256'hF960007000001C53EF66E557FFFFFFFFFFFFFFFFFEBFEEDFF23F4F7FFFFEFFFF;
defparam sdpb_inst_10.INIT_RAM_1A = 256'h7FE3043740000141FF7DE375FBFFFFFFFFFFFFFFFFF39F90FEEFF5F0FFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1B = 256'hA17F81081C000000FBFDEC3AAFEFFFFFFFFFFFFFFFFF78FB6FDBFFFF07FFFFFE;
defparam sdpb_inst_10.INIT_RAM_1C = 256'h3826FD0060E000021FF7FFE776FF7FFFFFFFFFFFFFFFF7BFE93E7B83E07FFFFF;
defparam sdpb_inst_10.INIT_RAM_1D = 256'hA5F92FE8111F800000FFFBFF18FBFFFFFFFFFFFFFFFFFFFCFFE47FBF3E07FFFD;
defparam sdpb_inst_10.INIT_RAM_1E = 256'hFB7A5BEF6050FC000023BBFFF37DFDFFFFFFFFFFFFFFFFFFC7DF93F8F3807FFF;
defparam sdpb_inst_10.INIT_RAM_1F = 256'hFD9E7EF1BB0883F0200279FFF80B16FFFFFFFFFFFFFFFFFFDE7CFEFF8F848FFF;
defparam sdpb_inst_10.INIT_RAM_20 = 256'hFFDF260AE5D8020FA0100FF7BBC4B9FFFFFFFFFFFFFFFBFFFF67AFFBF1FA88FF;
defparam sdpb_inst_10.INIT_RAM_21 = 256'hFFF9EBFF1AFEE8A13E6801EFFFBD2D36FFFFFFFFFFF7FBFFFFC83C3EFE9F509F;
defparam sdpb_inst_10.INIT_RAM_22 = 256'h7FFF343FFE4F760183FC800FCFFFFAA7FFFFFFFFFFFFBFFFDFFDFBE9EBC5E387;
defparam sdpb_inst_10.INIT_RAM_23 = 256'hE1FFF567FFFBD3A1240C73D4FFEFBE7B6FBFFFFFFFFFFFFEDDFFCFDFC7F1FE98;
defparam sdpb_inst_10.INIT_RAM_24 = 256'h951FFE2AFFFFD3FD40433DFD3FFFFFEFC17FFFFFFFFFDFFFFBE7FEFAFF147F99;
defparam sdpb_inst_10.INIT_RAM_25 = 256'h7C61FFEB8FFFFE8FE2007DFD7D6FF7ACA413FFFFFFFFFFDFFEDDDFFFAFB8CFA7;
defparam sdpb_inst_10.INIT_RAM_26 = 256'h8FEC0FFEF8FFFFF3BF501F7FD7FFF5FFBDA5FFFFFFFFFFFEFAEFFFFE399FE1FC;
defparam sdpb_inst_10.INIT_RAM_27 = 256'hE2FC01FFEF7FFFFF64FA83AFFFEFFAF7D64C7DFFFFFFFFFFF7678FFF07DE1FDF;
defparam sdpb_inst_10.INIT_RAM_28 = 256'h9E7F801FFE68FFFFF5CFDF5FFFFEFFFDFFEF7F7FFFFFFFFFFF9770D7E0FBFBF5;
defparam sdpb_inst_10.INIT_RAM_29 = 256'h5AFDBE03FFE3FFFFFF56FED7FFFFF7FF7FE4ECCFFFFFFFFFFFFFFE01FE07EFBF;
defparam sdpb_inst_10.INIT_RAM_2A = 256'hED6FC3C03FFF7F7FFFE74FEBFFFFFFFFFFDC81939FFFFFFFFFFFFF8017C07FFF;
defparam sdpb_inst_10.INIT_RAM_2B = 256'hE5FF7CFC07FFF3BBFFFCDEFEBFFFFFFFFFBFFD771FFFFFFFFFFFFDF82E7807F9;
defparam sdpb_inst_10.INIT_RAM_2C = 256'hEB3FDFC7007FFFB33FFF8DDFEBFFFFFFFFFFF3CC44B3FFFFFFFFFFFE90BE003F;
defparam sdpb_inst_10.INIT_RAM_2D = 256'h00007FFC400FFFFDBDFFF723FEA7FFFFFFFFFBABE012BFFFFFFFFFFFD81FE003;
defparam sdpb_inst_10.INIT_RAM_2E = 256'h800005F6B800FFFFE6EFF9EC7FE2FFFFFFEFFFFFF43C6FFFFFFFFFFFFDE7FE00;
defparam sdpb_inst_10.INIT_RAM_2F = 256'hFE00007F6E001FFFFEF67E6A8FFE7DFFFFFFFFF7BEC851FFFFFFFFFFFFBEF7F3;
defparam sdpb_inst_10.INIT_RAM_30 = 256'hEFF0000337C007FFFFF78EEAF1FFF57FFFFF8FFFDFB0E8AFFFFFFFFFFFFFC23E;
defparam sdpb_inst_10.INIT_RAM_31 = 256'hFEBE0000010000FFFFFF0F2AAB3FFF3BFFFFFEFFFFEE82D77FFFFFFFFFFF9C2F;
defparam sdpb_inst_10.INIT_RAM_32 = 256'hFFE8E000001C003FFFFFF9B3855FFFFBFFFFFEEFFFF9EEB85FFFFFFFFFFFFDC7;
defparam sdpb_inst_10.INIT_RAM_33 = 256'h07FC8E000007E047FFFFFFE506C7FFFF977FFFEAFFF7FDE003DFFFFFFFFFFF8D;
defparam sdpb_inst_10.INIT_RAM_34 = 256'h08FFBCE003BFFFFFFFFFFFFF931BFFFFFCB37FF7CFFFF313007FFFFFFFFFFFF8;
defparam sdpb_inst_10.INIT_RAM_35 = 256'hF007009E03FFFFFFFFFFFFFFFF003FFFFFE5BFDEE0FFFFF2D40BFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_36 = 256'hFE027FE9C07FFFFFFFFFFFFFFFFFFFFFF7FF33E23007FFF766F037FFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_37 = 256'hFFF038A0381FFFFFFFFFFFFFFFFFFFFFFDFFF8AD7A01FFFDFDC6BBFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_38 = 256'hFFFF03FC4703FFFFFFFFFFFFFFFFFFFFFFFFFFE332A047FFFF6E0FC7FFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_39 = 256'hFFFFF80CECE07FFFFFFFFFFFFFFFFFFFFFFEFFFF8738107FFFE6B6C9FFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3A = 256'hFFFFFFE074F807FFFFFFFFFFFFFFFFFFFFFFFD7FFE0C9249FF7F4EA01FFFFFFF;
defparam sdpb_inst_10.INIT_RAM_3B = 256'hFFFFFFFE80FE01DFFFFFFFFFFFFFFFFFFFFF3BFBFFFC150007E8FDBB86BFFFFF;
defparam sdpb_inst_10.INIT_RAM_3C = 256'hFFFFFFFFFC0000283FFFFFFFFFFFFFFFFFFFBF3FFFFFFCCA003D4FCB386FFFFF;
defparam sdpb_inst_10.INIT_RAM_3D = 256'hFFFFFFFFFFF8000301FFFFFFFFFFFFFFFFFFCD4FFFFFFFF60189EFEFFF0BEFFF;
defparam sdpb_inst_10.INIT_RAM_3E = 256'hFFFFFFFFFFFFE000BC1FFFFFFFFFFFFFFFFF853FFFFFFFFFB3140FFFBF7227FF;
defparam sdpb_inst_10.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFE207A9FFFFEFFFFFFFFFFF2C7FFFFFFFFFFD9042FB7B673BFF;

SDPB sdpb_inst_11 (
    .DO({sdpb_inst_11_dout_w[30:0],sdpb_inst_11_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_11.READ_MODE = 1'b1;
defparam sdpb_inst_11.BIT_WIDTH_0 = 1;
defparam sdpb_inst_11.BIT_WIDTH_1 = 1;
defparam sdpb_inst_11.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_11.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_11.RESET_MODE = "SYNC";
defparam sdpb_inst_11.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFA3FE5FFFEFFBFFFFFFC015FFFFFFFFFFFFEC884FF7FFE377;
defparam sdpb_inst_11.INIT_RAM_01 = 256'h2FFFFFFFFFFFFFFFFC0CF1FFFDFFFFFFFFA4FFFFFFFFFFFFFFFFA0583FFFDC67;
defparam sdpb_inst_11.INIT_RAM_02 = 256'hD9FFFFFFFFFFFFFFFF83CF9FFFBFFF7FFFE3FFFFFFFFFFFFFFFFFD2800FFFFFD;
defparam sdpb_inst_11.INIT_RAM_03 = 256'hDBBFFFFFFFFFFFFFFFF85C81FFFFFFFBFFF67FFFFFFFFFFDF7FFFFE934C7FFEF;
defparam sdpb_inst_11.INIT_RAM_04 = 256'hFBD7FFFFFFFFFFFFFFFF8F611FFFFFFFBFF3BFFFFFDFFF0FBF7FFFFF48103FFF;
defparam sdpb_inst_11.INIT_RAM_05 = 256'hFEF77FFFFFFFFFFFFFFFF8FE23FFFBFFF7F95FFFFEF972FC452FFFFFFA0101FF;
defparam sdpb_inst_11.INIT_RAM_06 = 256'h7FFFA7FFFFFFFFFFFFFFFF02E47FFFBFFF7E47FFFEEC7FFF7BBDFFFFFFD10C0F;
defparam sdpb_inst_11.INIT_RAM_07 = 256'h03FFDFFFFFFFFFFFFFFFFFE19E9FFFFFFFCFC9FFFF2DFFFFBCFF30DFFFFE8208;
defparam sdpb_inst_11.INIT_RAM_08 = 256'h821FFFD7FFFFFFFFFFFFFFFE77D1FFFFDFF9EA7FFFBEFFFFF4E6DFC69FFFF402;
defparam sdpb_inst_11.INIT_RAM_09 = 256'h0081FFF3FFFFFFFFFFFFFFFFC7FA3FFFFFFF791FFFEE7FFFFF84FE9807DFFFA0;
defparam sdpb_inst_11.INIT_RAM_0A = 256'hE8308FFFFFFFFFFFFFFFFFFFFC3647FFFFFFCF17FFFB9FFFFFF17FFF9C7B7FFD;
defparam sdpb_inst_11.INIT_RAM_0B = 256'hFF40203FFFFFFFFFFFFFFFFFFF8A58FFFFFF378CFFFFAFFFFFFC1FFFFF697FFF;
defparam sdpb_inst_11.INIT_RAM_0C = 256'hFFFA0433FFF7FFFFFFFFFFFFFFF31B9FFFFFFCF7BFFF33FFFFFF85FFFFFD437F;
defparam sdpb_inst_11.INIT_RAM_0D = 256'hFFFFF00C1FFF7FFFFFFFFFFFFFFE6F53FFFFFFFFF7FFD8FFFFFFF07FFFFFEE1F;
defparam sdpb_inst_11.INIT_RAM_0E = 256'h8FFFFF830CFFFFFFFFFFFFFFFFFFC7A23FFFFFFFCCFFF57FFFFFFF87FFFFFFA1;
defparam sdpb_inst_11.INIT_RAM_0F = 256'hE87FFFFC030BFFCFFFFFFFFFFFFFF832C7FFFFFFFD1FFEFFFFFFFFF07FFFFFFF;
defparam sdpb_inst_11.INIT_RAM_10 = 256'hFFCBFFFFE0831FFFFFFFFFFFFFFFFF8A747FFFFFFF83FFB7FFFFFFFF07FFFFFF;
defparam sdpb_inst_11.INIT_RAM_11 = 256'hFFF61FFFFF00C2FFFFFFFFFFFFFFFFF1DC8FFFFFFFF17FEFFFFFFFFFF47FFFFF;
defparam sdpb_inst_11.INIT_RAM_12 = 256'hFFFFB9FFFFF02407FFFFFFFFFFFFFFFC6DB0FFFFFFFE6FFFFFFFFFFFFE67FFFF;
defparam sdpb_inst_11.INIT_RAM_13 = 256'hFFFFFB8FFFFFC410BFFFFFFFFFFFFFFF8F9D1FFFFFFFF5FFB3FFFFFFFFEE7FFF;
defparam sdpb_inst_11.INIT_RAM_14 = 256'hFFFFFFD8FFFFFC0021FFFFFFFFFFFFFFF0DA21FFFFFFFA9FF27FFFFFFFFF63FF;
defparam sdpb_inst_11.INIT_RAM_15 = 256'hFFFFFFFFCFFFFFE80C2FFFFFFFFFFFFFFC09CE3FFFFFFF83FE47FFFFFFFFF73F;
defparam sdpb_inst_11.INIT_RAM_16 = 256'h3FFFFFFFE87FFFFF02207FFFFFFFFFFFFF81C7C3FFFFFFF13FCE7FFFFFFFFFBD;
defparam sdpb_inst_11.INIT_RAM_17 = 256'hFFFFFFFFFE97FFFFF84101FFFFFFFFFFFFE07AE87FFFFFFEE7F9CFFFFFFFFFF9;
defparam sdpb_inst_11.INIT_RAM_18 = 256'hFD67FFFFFFE17FFFFFC0580FFFFFFFFFFFF037D987FFFFFFDCFF90FFFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_19 = 256'hFFE77FFFFFFE0FFFFFFE9430FFFFFFFFFFFCE6F7D07FFFFFF81FF29FFFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1A = 256'hFFFF7EFFFFFFD8FFFFFFF00057FFFFFFFFFEEFDC3B0FFFFFFF89FE51FFFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1B = 256'hFFFFF9CFFFFFFC1FFFFFFFA4803FFFFFFFFFFC5EF4A0FFFFFFF01FCC3FFFFFFF;
defparam sdpb_inst_11.INIT_RAM_1C = 256'hFFFFFFF77FFFFF81FFFFFFFD0400FFFFFFFFF61F4DF30FFFFFFF67F8A3FFFFFF;
defparam sdpb_inst_11.INIT_RAM_1D = 256'hFFFFFFFE5AFFFFB83FFFFFFFE10087FFFFFFFE83FF92307FFFFFEE7F047FFFFF;
defparam sdpb_inst_11.INIT_RAM_1E = 256'hFFFFFFFFF1FFFFD487FFFFFFFE00003FFFFFFFC836930187FFFFFE4FF1C7FFFF;
defparam sdpb_inst_11.INIT_RAM_1F = 256'hFFFFFFFFFF97FFBEFEFFFFFFFFF01801FFFFFFF5077CE07C3FFFFFD4FE087FFF;
defparam sdpb_inst_11.INIT_RAM_20 = 256'hFFFFFFFFFF3E5DBFFF1FFFFFFFFFC0006FFFFFFF10FFEE0643FFFFF89FC30FFF;
defparam sdpb_inst_11.INIT_RAM_21 = 256'hFFFFFFFFA00931C7FF8FFFFFFFFFFC80DC7FFFFFF11FFDC0163FFFFF81F8507F;
defparam sdpb_inst_11.INIT_RAM_22 = 256'hFFFFFFFFC00002806D87FFFFFFFFFFE08207FFFFFE3FFF1E01E1FFFFFB1F860F;
defparam sdpb_inst_11.INIT_RAM_23 = 256'h0FFFFFFFC00020090007FFFFFFFFFFFF30C03FFFFFC3F7EEC06A1FFFFF03F060;
defparam sdpb_inst_11.INIT_RAM_24 = 256'hC07FFFFF4000DD00A0FFFFFFFFFFFFFFF93403FFFFFC67FB8C07C1FFFFF53E0E;
defparam sdpb_inst_11.INIT_RAM_25 = 256'h0C07FFFFCC0019000101FFFFFFFFFFFFFFDC001FFFFF80FCEB00A407FFFF6700;
defparam sdpb_inst_11.INIT_RAM_26 = 256'h00403FFFFE00066F40040FFFFFFFFFFFFFFEC003FFFFE0DFEAE01740FFFFE650;
defparam sdpb_inst_11.INIT_RAM_27 = 256'h001C09FFFF8001DFFE1058FFFFFFFFFFFFFFF5003FFFFD0697FE06C807FFFF24;
defparam sdpb_inst_11.INIT_RAM_28 = 256'h08018017FFFC0018BFE70103FFFFFFFFFFFFFFC817FFFF23227F007900FFFFC8;
defparam sdpb_inst_11.INIT_RAM_29 = 256'h84401809FFDDC00712FFDC0E0FFFFFFFFFFFFFFF25FFFFDC23881016301FFFF8;
defparam sdpb_inst_11.INIT_RAM_2A = 256'hF000018009EF5000E35FFF38EB7FFFFFFFFFFFFFFFFFFFFBDE302002C601FFFF;
defparam sdpb_inst_11.INIT_RAM_2B = 256'hBE1400280078E0001EFFFFDBE32BFFFFFFFFFFFFFFFFFFFE7BA781801DC00BFF;
defparam sdpb_inst_11.INIT_RAM_2C = 256'hFCC0C000800EC90003DDFFFBE7BC8FFFFFFFFFFFFFFFFFFFCFF1357B47B801FF;
defparam sdpb_inst_11.INIT_RAM_2D = 256'h796C1400380044020078D7FFFDBBDA3FFFFFFFFFFFFFFFFBD1FCFDCEF8E58011;
defparam sdpb_inst_11.INIT_RAM_2E = 256'h10E8824003800108000714FFF7BFCADEFFFFFFFFFFFFFFFFFE1FAFA749AF5000;
defparam sdpb_inst_11.INIT_RAM_2F = 256'h00000004007000000000F3215EFFDFBA47FFFFFFFFFFFFFFFBC3793C7D88F300;
defparam sdpb_inst_11.INIT_RAM_30 = 256'h000002004001000000000EBFDFDF7BDEFD1FFFFFFFFFFFFFFEC83E7004287FB0;
defparam sdpb_inst_11.INIT_RAM_31 = 256'hA000000028007000000000EB7F7DEFFFFB60FFFFFFFFFFFFFFF90FAF031503FB;
defparam sdpb_inst_11.INIT_RAM_32 = 256'hBA00000001C007000000001D6FF7BFF77FF9037BFFFFFFFFFFFF407C6007743F;
defparam sdpb_inst_11.INIT_RAM_33 = 256'h0BA000000008003000000001DCF777DEFFFFA6059BFF7FFFFFFFF40FC1707903;
defparam sdpb_inst_11.INIT_RAM_34 = 256'h006A000000038003000000001D76A3BFFF3BFFCC107FDFFFFFFFF640FD000380;
defparam sdpb_inst_11.INIT_RAM_35 = 256'h000CE00000001801A000000001D7A68CBDE287FCB30FFFEFFFFFF5E00B800008;
defparam sdpb_inst_11.INIT_RAM_36 = 256'h00007400000005800E000000001D398133FE000FFDB0017D9FFFBEFE40FC8000;
defparam sdpb_inst_11.INIT_RAM_37 = 256'h0000DDC000000078036000000001D3E6024382000EFFC015FFFFFF2F7003C000;
defparam sdpb_inst_11.INIT_RAM_38 = 256'h000019E8000000038036000000000C9F5804080000FCC8003FC5FFF328007C00;
defparam sdpb_inst_11.INIT_RAM_39 = 256'h90000731800000003806C000000000E57590116400077B94012F1FFD7E0803E0;
defparam sdpb_inst_11.INIT_RAM_3A = 256'hBF1800EF7000000001806C000000000F689AF1590000D03FD0021A458100003F;
defparam sdpb_inst_11.INIT_RAM_3B = 256'h0E3F02304E00000001D80EC0000000007B233081E0000EC06480000080000001;
defparam sdpb_inst_11.INIT_RAM_3C = 256'h0072F9D8DCE00000003D80F80000000007D87B591D8000BFFEF40004B4018000;
defparam sdpb_inst_11.INIT_RAM_3D = 256'h0001C818BE5C00000007FC3F80000000003E56EF4CC0003DFFBF200000000800;
defparam sdpb_inst_11.INIT_RAM_3E = 256'h00000794255300000000CEFF980000000001F36FF76F68015FFB088000000000;
defparam sdpb_inst_11.INIT_RAM_3F = 256'h0000001E34C9E00000000CDFFD80000000000FCD3FD7F1800BFFF3F400000000;

SDPB sdpb_inst_12 (
    .DO({sdpb_inst_12_dout_w[30:0],sdpb_inst_12_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_12.READ_MODE = 1'b1;
defparam sdpb_inst_12.BIT_WIDTH_0 = 1;
defparam sdpb_inst_12.BIT_WIDTH_1 = 1;
defparam sdpb_inst_12.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_12.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_12.RESET_MODE = "SYNC";
defparam sdpb_inst_12.INIT_RAM_00 = 256'hDFFFFFFFFFFFFFFFFF20100000001BFFFFFFFFFFFF7FFDFDFFFFFFFFFFFFFFFE;
defparam sdpb_inst_12.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFE2000C000009AFFFFFFFFFFFFF6FE3AFFFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFD000300000002BF7FFFFF7B860C03C5DFFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFA080080400000637EFFFA82028004861CFB7FFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFF8400300100004010F05C9000000011C4407FFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFE0002001F000100772B00B200000115401FFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFEF0000FC03080000473A1864000000003806EFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFF82071F1F030040DBF9A0600000000906E5A7FFFFF;
defparam sdpb_inst_12.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE800007F800801C17FA50000000000100777FFFFF;
defparam sdpb_inst_12.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC03001F000FFEE9FF7B06004000800800BDFFFF;
defparam sdpb_inst_12.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE400003FC01CFFFB77FB480540B0000417BF6FB;
defparam sdpb_inst_12.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE827003DF0703FFFFFFF8000002350002FEDAF;
defparam sdpb_inst_12.INIT_RAM_0C = 256'h71FEFF9FFFFFFFFFFFFFFFFFFFFF223E1E07EF00FFFFFDF0000000B500006EED;
defparam sdpb_inst_12.INIT_RAM_0D = 256'hEFFFFFFFFFFFFFFFFFFFFFFFFFFF5C01F5C01FC003FFFFFE00007C100081046F;
defparam sdpb_inst_12.INIT_RAM_0E = 256'h6FDFFFFFFFFFFFFFFFFFFFFFFFFFFFF007F8007C00EFFFFFE0103E1C28E8004F;
defparam sdpb_inst_12.INIT_RAM_0F = 256'hA7DBFF3FFFFFFFFFFFFFFFFFFFFFFFAE003F001EF80EFFFFFA000E0A7000B023;
defparam sdpb_inst_12.INIT_RAM_10 = 256'h00CE1EF29FFFFBFFFFFFFFFFFFFFFFFFC007DC0387C7CFFFFF000387A7000100;
defparam sdpb_inst_12.INIT_RAM_11 = 256'h00077FFFFBFFFDFFFFFFFFFFFFFFFFFFFE00E0F8F81F61FFFFF44030D81A0000;
defparam sdpb_inst_12.INIT_RAM_12 = 256'h00000A7FF7EFEFFDFBFFFFFFFFFFFFFFFF983E03BE007E1FFFFF200F20107000;
defparam sdpb_inst_12.INIT_RAM_13 = 256'h00000003BFDBFF97FFFFFFFFFFFFFFFFFFEF6F800DC00300FFFFF006F8080380;
defparam sdpb_inst_12.INIT_RAM_14 = 256'hE00188017EFFDFF7FFFFFFFFFFFFFFFFFFFFBBF003FE00E81FFFFD842FCA001C;
defparam sdpb_inst_12.INIT_RAM_15 = 256'h8E001F00003F6DFEFFFFDFFFFFFFFFFFFFFFFFE6003FF80E00FFFFF000FE003B;
defparam sdpb_inst_12.INIT_RAM_16 = 256'h847803048C17BFFE3C9FF7FFFFFFFFFFFFFFFFDF3C0B8BE7084FFFFF8007F81F;
defparam sdpb_inst_12.INIT_RAM_17 = 256'h810B800000DFBFFFF77DFFFFFFFFFFFFFFFFFFFFFAE1F00F6083FFFFFE017F84;
defparam sdpb_inst_12.INIT_RAM_18 = 256'hBC881E00000007FBC7A38FF7FFFFFFFFFFFFFFFFEF1BDC00BC084FFFFF740FF0;
defparam sdpb_inst_12.INIT_RAM_19 = 256'hFE21287000001C53EF66E557FFFFFFFFFFFFFFFFFF3BFFA00F0000FFFFFEFFFF;
defparam sdpb_inst_12.INIT_RAM_1A = 256'hFFF90C3740000141FF7DE375FBFFFFFFFFFFFFFFFFF5DFFF0158080FFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1B = 256'h5F7FD1003C000000FBFDEC3AAFEFFFFFFFFFFFFFFFFF70FCF0388100FFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_1C = 256'h519BFE8021E000021FF7FFE776FF7FFFFFFFFFFFFFFFFF9FCBC708481FFFFFFE;
defparam sdpb_inst_12.INIT_RAM_1D = 256'hD80093F41947800000FFFBFF18FBFFFFFFFFFFFFFFFFFFFE7CEFC08282FFFFFE;
defparam sdpb_inst_12.INIT_RAM_1E = 256'hF08C201FA050BC000023BBFFF37DFDFFFFFFFFFFFFFFFFFFCDCFBC00487FFFFF;
defparam sdpb_inst_12.INIT_RAM_1F = 256'hFE6603437D0841F0200279FFF80B16FFFFFFFFFFFFFFFFFFFE65FF0080377FFF;
defparam sdpb_inst_12.INIT_RAM_20 = 256'hFFF09FF081E8128FA0100FF7BBC4B9FFFFFFFFFFFFFFF3FFFC77D7E4000277FF;
defparam sdpb_inst_12.INIT_RAM_21 = 256'hFFFE17FFE85F40A17E6801EFFFBD2D36FFFFFFFFFFFFFFDFFFC07D3F4000CF7F;
defparam sdpb_inst_12.INIT_RAM_22 = 256'hFFFFC8FFFFB07A1001FC800FCFFFFAA7FFFFFFFFFFFFBFBFFDFF83E7E04C127F;
defparam sdpb_inst_12.INIT_RAM_23 = 256'h5FFFFA3FFFFC0FC0051FF3D4FFEFBE7B6FBFFFFFFFFFFFBBFDFFEE1F77084286;
defparam sdpb_inst_12.INIT_RAM_24 = 256'h0AFFFFD1FFFFE89E0042C27D3FFFFFEFC17FFFFFFFFFDFFBEFFFFFF8F7FA0440;
defparam sdpb_inst_12.INIT_RAM_25 = 256'h049FFFF47FFFFF61F8208202FD6FF7ACA413FFFFFFFFFFDFFFFDFFFFA3BB1014;
defparam sdpb_inst_12.INIT_RAM_26 = 256'h1053FFFF03FFFFF85F8000006BFFF5FFBDA5FFFFFFFFFFFEFFEF9FFFF9F3FC04;
defparam sdpb_inst_12.INIT_RAM_27 = 256'h130BFFFFF49FFFFF81FC0C50000FFAF7D64C7DFFFFFFFFFDFF7FFF7FF8CFDFA0;
defparam sdpb_inst_12.INIT_RAM_28 = 256'hC2B07FFFFFD1FFFFFA3FEAA000017FFDFFEF7F7FFFFFFFFFFFFFFFF7FF03FDF2;
defparam sdpb_inst_12.INIT_RAM_29 = 256'h9D5161FFFFF80FFFFFA9FF5800000FFF7FE4ECCFFFFFFFFFFFEFFFFFFFF81F8F;
defparam sdpb_inst_12.INIT_RAM_2A = 256'hCC18083FFFFFB0FFFFF81FF30000003FFFDC81939FFFFFFFFFFFFFFFF7FF807C;
defparam sdpb_inst_12.INIT_RAM_2B = 256'h16F00203FFFFFC0FFFFFA1FF20000003FFBFFD771FFFFFFFFFFFFDFFD13FF805;
defparam sdpb_inst_12.INIT_RAM_2C = 256'h14EFE038FFFFFFD5BFFFE03FF30000009FFFF3CC44B3FFFFFFFFFFFE7F01FFC0;
defparam sdpb_inst_12.INIT_RAM_2D = 256'hFFFF7C07BFFFFFFEC7FFFAD7FF28000000FFFBABE012BFFFFFFFFFFFC7E01FFC;
defparam sdpb_inst_12.INIT_RAM_2E = 256'h7FFFF9E9C7FFFFFFF01FFE02FFFA0000000FFFFFF43C6FFFFFFFFFFFFE1800FF;
defparam sdpb_inst_12.INIT_RAM_2F = 256'h81FFFF8EA1FFFFFFFF4CFF845FFFA2000000FFF7BEC851FFFFFFFFFFFFC10814;
defparam sdpb_inst_12.INIT_RAM_30 = 256'h180FFFFCA03FFFFFFFFA41140BFFF80000007FFFDFB0E8AFFFFFFFFFFFF83DC1;
defparam sdpb_inst_12.INIT_RAM_31 = 256'h0181FFFFFE7FFFFFFFFFC0C41AFFFFD0000001FFFFEE82D77FFFFFFFFFFFE3D0;
defparam sdpb_inst_12.INIT_RAM_32 = 256'h00181FFFFFFFFFFFFFFFFECC0B3FFFFCA020017FFFF9EEB85FFFFFFFFFFFFC38;
defparam sdpb_inst_12.INIT_RAM_33 = 256'hF80381FFFFFFFFFFFFFFFFF8CBDFFFFFE500001DFFF7FDE003DFFFFFFFFFFFD3;
defparam sdpb_inst_12.INIT_RAM_34 = 256'hFF003C1FFFFFFFFFFFFFFFFFE017FFFFFF2000003FFFF313007FFFFFFFFFFFFE;
defparam sdpb_inst_12.INIT_RAM_35 = 256'hFFB8FF81FFFFFFFFFFFFFFFFFFFFBFFFFFF9002005FFFFF2D40BFFFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_36 = 256'hFFFCBF983FFFFFFFFFFFFFFFFFFFFFFFF7FFC51D080FFFF766F037FFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_37 = 256'hFFFFC0FB07FFFFFFFFFFFFFFFFFFFFFFFDFFFF3182017FFDFDC6BBFFFFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_38 = 256'hFFFFFC3B60FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC392063FFFF6E0FC7FFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_39 = 256'hFFFFFFF0F41FFFFFFFFFFFFFFFFFFFFFFFFEFFFFF800105FFFE6B6C9FFFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3A = 256'hFFFFFFFF8407FFFFFFFFFFFFFFFFFFFFFFFFFD7FFFF18818FF7F4EA01FFFFFFF;
defparam sdpb_inst_12.INIT_RAM_3B = 256'hFFFFFFFFFF01FFFFFFFFFFFFFFFFFFFFFFFFA7FBFFFFEC040FE8FDBB86BFFFFF;
defparam sdpb_inst_12.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFFFFFF42047D4FCB386FFFFF;
defparam sdpb_inst_12.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFE27FFFFFFFFA040BEFEFFF0BEFFF;
defparam sdpb_inst_12.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFF23FFFFFFFFFFFFFFFFFFE0FFFFFFFFFFD1051FFFBF7227FF;
defparam sdpb_inst_12.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFCF7FFFFFFFFFFFFFFFE85FFFFFFFFFFFE8122FB7B673BFF;

SDPB sdpb_inst_13 (
    .DO({sdpb_inst_13_dout_w[30:0],sdpb_inst_13_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_13.READ_MODE = 1'b1;
defparam sdpb_inst_13.BIT_WIDTH_0 = 1;
defparam sdpb_inst_13.BIT_WIDTH_1 = 1;
defparam sdpb_inst_13.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_13.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_13.RESET_MODE = "SYNC";
defparam sdpb_inst_13.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFC9F3FFFFFFFFFFFFFF033FFFFFFFFFFFFF44147F7FFE377;
defparam sdpb_inst_13.INIT_RAM_01 = 256'h2FFFFFFFFFFFFFFFFFFB07FFFFFFEFFFFFC1FFFFFFFFFFFFFFFFE0083FFFDC67;
defparam sdpb_inst_13.INIT_RAM_02 = 256'hD9FFFFFFFFFFFFFFFFFB197FFFFFFF7FFFE5FFFFFFFFFFFFFFFFFF1040FFFFFD;
defparam sdpb_inst_13.INIT_RAM_03 = 256'hDBBFFFFFFFFFFFFFFFFFFE6FFFFBFFFFFFE3FFFFFFFFFFFEAFFFFFF820C7FFEF;
defparam sdpb_inst_13.INIT_RAM_04 = 256'hFBD7FFFFFFFFFFFFFFFFF07CFFFFBFFFFFF97FFFFFF800F0007FFFFFC4203FFF;
defparam sdpb_inst_13.INIT_RAM_05 = 256'hFEF77FFFFFFFFFFFFFFFFFE99FFFFFFFF7FC3FFFFF030D00071FFFFFFE0C21FF;
defparam sdpb_inst_13.INIT_RAM_06 = 256'h7FFFA7FFFFFFFFFFFFFFFFED13FFFFFFFFFE5FFFFF9BFFFF84423FFFFFF1000F;
defparam sdpb_inst_13.INIT_RAM_07 = 256'h03FFDFFFFFFFFFFFFFFFFFFDE27FFFFFFFDFC7FFFF8BFFFFC300CF5FFFFF8140;
defparam sdpb_inst_13.INIT_RAM_08 = 256'h501FFFD7FFFFFFFFFFFFFFFF8E4FFFFFFFFBE1FFFFC5FFFFFB10003B9FFFFC01;
defparam sdpb_inst_13.INIT_RAM_09 = 256'h0041FFF3FFFFFFFFFFFFFFFFFC49FFFFFFFFFD7FFFF8FFFFFF7BFF63FFDFFFE0;
defparam sdpb_inst_13.INIT_RAM_0A = 256'hF8140FFFFFFFFFFFFFFFFFFFFFC33FFFFFFFDF0FFFFCFFFFFFEEFFFFE3FB7FFF;
defparam sdpb_inst_13.INIT_RAM_0B = 256'hFFC0107FFFFFFFFFFFFFFFFFFFEDB7FFFFFFB3E3FFFE1FFFFFFFFFFFFF967FFF;
defparam sdpb_inst_13.INIT_RAM_0C = 256'hFFFE0511FFF7FFFFFFFFFFFFFFFEF67FFFFFFFFC7FFFDFFFFFFFFBFFFFFEBF7F;
defparam sdpb_inst_13.INIT_RAM_0D = 256'hFFFFF0000FFF7FFFFFFFFFFFFFFF924FFFFFFFFF8FFFE3FFFFFFFFFFFFFFF1FF;
defparam sdpb_inst_13.INIT_RAM_0E = 256'h7FFFFF81447FFFFFFFFFFFFFFFFFF859FFFFFFFFE3FFFAFFFFFFFFFFFFFFFFDF;
defparam sdpb_inst_13.INIT_RAM_0F = 256'hF7FFFFFC000BFFCFFFFFFFFFFFFFFFEDBFFFFFFFFE7FFF3FFFFFFFFFFFFFFFFE;
defparam sdpb_inst_13.INIT_RAM_10 = 256'hFF37FFFFE0511FFFFFFFFFFFFFFFFFE513FFFFFFFFCFFFDFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_11 = 256'hFFF9FFFFFF0002FFFFFFFFFFFFFFFFFE167FFFFFFFF8FFF1FFFFFFFFFBFFFFFF;
defparam sdpb_inst_13.INIT_RAM_12 = 256'hFFFFC7FFFFF010C7FFFFFFFFFFFFFFFF926FFFFFFFFF5FFE3FFFFFFFFF9FFFFF;
defparam sdpb_inst_13.INIT_RAM_13 = 256'hFFFFFC7FFFFFC420BFFFFFFFFFFFFFFFF064FFFFFFFFEBFFC7FFFFFFFFF1FFFF;
defparam sdpb_inst_13.INIT_RAM_14 = 256'hFFFFFFE7FFFFFC0D31FFFFFFFFFFFFFFFF389FFFFFFFFC7FFCFFFFFFFFFF9FFF;
defparam sdpb_inst_13.INIT_RAM_15 = 256'hFFFFFFFE3FFFFFE9082FFFFFFFFFFFFFFFF3B9FFFFFFFFCFFF9FFFFFFFFFF8FF;
defparam sdpb_inst_13.INIT_RAM_16 = 256'hDFFFFFFFF7FFFFFF03647FFFFFFFFFFFFFFD393FFFFFFFF8FFF5FFFFFFFFFFC3;
defparam sdpb_inst_13.INIT_RAM_17 = 256'hC1FFFFFFFF7FFFFFF80003FFFFFFFFFFFFFFC627FFFFFFFF5FFF3FFFFFFFFFFE;
defparam sdpb_inst_13.INIT_RAM_18 = 256'hFE1FFFFFFFFFFFFFFFC0110FFFFFFFFFFFFFC08C7FFFFFFFE3FFE7FFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_19 = 256'hFFF8FFFFFFFFFFFFFFFE8470FFFFFFFFFFFF102C4FFFFFFFFE7FFC7FFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1A = 256'hFFFF81FFFFFFE7FFFFFFF01053FFFFFFFFFF1007C8FFFFFFFFF7FFEFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1B = 256'hFFFFFE3FFFFFFFFFFFFFFFA1821FFFFFFFFFC3A5819FFFFFFFFCFFF1FFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1C = 256'hFFFFFFE0BFFFFFFFFFFFFFFD0404FFFFFFFFFDE02350FFFFFFFFFFFF1FFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1D = 256'hFFFFFFFF85FFFFC7FFFFFFFFE16007FFFFFFFF7C024D0FFFFFFFF1FFEBFFFFFF;
defparam sdpb_inst_13.INIT_RAM_1E = 256'hFFFFFFFFFC007FEB7FFFFFFFFF00113FFFFFFFF7C978F87FFFFFFF7FFE3FFFFF;
defparam sdpb_inst_13.INIT_RAM_1F = 256'hFFFFFFFFFFE4004101FFFFFFFFF81001FFFFFFFEF8E7DFA3FFFFFFE3FFE7FFFF;
defparam sdpb_inst_13.INIT_RAM_20 = 256'hFFFFFFFFFFFF840000FFFFFFFFFFC0046FFFFFFFEF3C19FA3FFFFFFEFFFCFFFF;
defparam sdpb_inst_13.INIT_RAM_21 = 256'hFFFFFFFFFFEEFE04007FFFFFFFFFFE80D47FFFFFFCE703BFC1FFFFFFE7FF8FFF;
defparam sdpb_inst_13.INIT_RAM_22 = 256'hFFFFFFFFFFFDFDFF807FFFFFFFFFFFF00107FFFFFFC060FDFD9FFFFFFEFFF9FF;
defparam sdpb_inst_13.INIT_RAM_23 = 256'hFFFFFFFFFFFF7FF7FFFFFFFFFFFFFFFFB0403FFFFFFC0610FFB9FFFFFFCFFF5F;
defparam sdpb_inst_13.INIT_RAM_24 = 256'h3FFFFFFFFFFF33FFDFFFFFFFFFFFFFFFFD1403FFFFFF98E47BF8BFFFFFF8FFF1;
defparam sdpb_inst_13.INIT_RAM_25 = 256'hEBFFFFFFFFFFE6FFFFFFFFFFFFFFFFFFFFEC003FFFFFFA861F7F53FFFFFFDFFF;
defparam sdpb_inst_13.INIT_RAM_26 = 256'hFE3FFFFFFFFFF89FFFFEFFFFFFFFFFFFFFFF4003FFFFFEE07AEFE13FFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_27 = 256'hFFE3FFFFFFFFFE03FDFFB7FFFFFFFFFFFFFFF9007FFFFE8369FDFC67FFFFFF9F;
defparam sdpb_inst_13.INIT_RAM_28 = 256'h3FFE7FFFFFFFFFE37FF7FEFFFFFFFFFFFFFFFFE00FFFFFC27D80FFACFFFFFFF3;
defparam sdpb_inst_13.INIT_RAM_29 = 256'hF7FFE7FFFFFFFFF84FFE5FF7FFFFFFFFFFFFFFFFC3FFFFE05877EFE08FFFFFFF;
defparam sdpb_inst_13.INIT_RAM_2A = 256'hFF3FFE7FFFFFFFFF06FFC13F2FFFFFFFFFFFFFFFFFFFFFFC538FDFFC11FFFFFF;
defparam sdpb_inst_13.INIT_RAM_2B = 256'hFFE3FFD7FFFFFFFFE01FF801FCB7FFFFFFFFFFFFFFFFFFFF845C7E7FC33FFFFF;
defparam sdpb_inst_13.INIT_RAM_2C = 256'hFFFE3FFF7FFFFFFFFC0BFF800FC0FFFFFFFFFFFFFFFFFFFFF00E8A94B867FFFF;
defparam sdpb_inst_13.INIT_RAM_2D = 256'hFFFFEBFFC7FFFFFFFF81BFF0003E3DFFFFFFFFFFFFFFFFFFFE030431070C7FFF;
defparam sdpb_inst_13.INIT_RAM_2E = 256'hFFFFFC3FFC7FFFFFFFF83BFE0001F9E7FFFFFFFFFFFFFFFFFFC05050B610CFFF;
defparam sdpb_inst_13.INIT_RAM_2F = 256'hFFFFFFE3FF8FFFFFFFFF05F9600007E5FFFFFFFFFFFFFFFFFFF814E3667708FF;
defparam sdpb_inst_13.INIT_RAM_30 = 256'hFFFFFFFE3FFCFFFFFFFFF0FFF800003FC7FFFFFFFFFFFFFFFFFF85887FD7C08F;
defparam sdpb_inst_13.INIT_RAM_31 = 256'h9FFFFFFFC7FF8FFFFFFFFF0FFF800007FF1FFFFFFFFFFFFFFFFFF04003FAFC08;
defparam sdpb_inst_13.INIT_RAM_32 = 256'h09FFFFFFFC3FF8FFFFFFFFE17FFC00007FF857FFFFFFFFFFFFFFFF0300068BC0;
defparam sdpb_inst_13.INIT_RAM_33 = 256'hF09FFFFFFFC7FF4FFFFFFFFE17F7F8000FFFE3FFFFFFFFFFFFFFFFF83F7002FE;
defparam sdpb_inst_13.INIT_RAM_34 = 256'hFF59FFFFFFFE7FF8FFFFFFFFE18EB3B0013BFF83FFFFFFFFFFFFFFFF82FFFC7F;
defparam sdpb_inst_13.INIT_RAM_35 = 256'hFFF39FFFFFFFC7FE1FFFFFFFFE18668C800287FF8EFFFFFFFFFFFFFFF47FFFFF;
defparam sdpb_inst_13.INIT_RAM_36 = 256'hFFFF93FFFFFFF87FE1FFFFFFFFE1C7FF3202100FFF0FFFFFFFFFFFFFFF037FFF;
defparam sdpb_inst_13.INIT_RAM_37 = 256'hFFFFE33FFFFFFFA7FC1FFFFFFFFE1C1FFE4402000E18FFFFFFFFFFFFFFF83FFF;
defparam sdpb_inst_13.INIT_RAM_38 = 256'hFFFFDD27FFFFFFF87FC1FFFFFFFFF0E0FFFD180000E0177FFFFFFFFFFFFF83FF;
defparam sdpb_inst_13.INIT_RAM_39 = 256'h77FFFD047FFFFFFF87FB3FFFFFFFFF068BDFF7640006802BFFFFFFFFFFFFFC1F;
defparam sdpb_inst_13.INIT_RAM_3A = 256'h00DFFF41CFFFFFFFF07F83FFFFFFFFF0786FFF798000CFC0EFFFFFFFFFFFFFCC;
defparam sdpb_inst_13.INIT_RAM_3B = 256'hF045C3B099FFFFFFFF07F03FFFFFFFFF83FDDE01E0000DFF8F3FFFFFFFFFFFFE;
defparam sdpb_inst_13.INIT_RAM_3C = 256'hFF80073CA21FFFFFFFC07F47FFFFFFFFF81C96F0078000DFFCFBFFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3D = 256'hFFFE09E708C3FFFFFFF823C27FFFFFFFFFC06419403E003BFFCFDFFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3E = 256'hFFFFF81456B0FFFFFFFF020087FFFFFFFFFE03A82E103801BFFC7FFFFFFFFFFF;
defparam sdpb_inst_13.INIT_RAM_3F = 256'hFFFFFFE038381FFFFFFFF040007FFFFFFFFFF00E20B010C007FF87FBFFFFFFFF;

SDPB sdpb_inst_14 (
    .DO({sdpb_inst_14_dout_w[29:0],sdpb_inst_14_dout[5:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[15],ada[14],ada[13]}),
    .BLKSELB({adb[15],adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_14.READ_MODE = 1'b1;
defparam sdpb_inst_14.BIT_WIDTH_0 = 2;
defparam sdpb_inst_14.BIT_WIDTH_1 = 2;
defparam sdpb_inst_14.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_14.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_14.RESET_MODE = "SYNC";
defparam sdpb_inst_14.INIT_RAM_00 = 256'hAAAAAAAAAAAA95550E96555ADD5C1532003D6BFFFF952FFBAAAAAAAAAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_01 = 256'hAAAAAAAAAAAAAAAA95540000556AAAAAAAAAAAAAAAAA55715550115AAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_02 = 256'hAAAAAAAAAAAAAAA95540E914556DA0555273F5AFFFFE552FFBEAAAAAAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_03 = 256'hAAAAAAAAAAAAAAAAAAA955555556AAAAAAAAAAAAAAAAA575715550616AAAAAAA;
defparam sdpb_inst_14.INIT_RAM_04 = 256'hAAAAAAAAAAAAAAAAAA55543E454556D041452FD6ABFFFE55EBFBFBAAAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_05 = 256'hAAAAAAAAAAAAAAAAAAAAAAAA659AAAAAAAAAAAAAAAAAAAA951C55548716AAAAA;
defparam sdpb_inst_14.INIT_RAM_06 = 256'hAAAAAAAAAAAAAAAAAAAAA55543E454AA790050AF5AABFFFD14BFA8CEAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_07 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55E055540B16AAA;
defparam sdpb_inst_14.INIT_RAM_08 = 256'hAAAAAAAAAAAAAAAAAAAAAAA555543E556A971105571AABFFF914BFF97FAAAAAA;
defparam sdpb_inst_14.INIT_RAM_09 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA955555544056A;
defparam sdpb_inst_14.INIT_RAM_0A = 256'h6AAAAAAAAAAAAAAAAAAAAAAAA9555543E432A970414846AFFFF855FFFEA1AAAA;
defparam sdpb_inst_14.INIT_RAM_0B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5556554085;
defparam sdpb_inst_14.INIT_RAM_0C = 256'hC5AAAAAAAAAAAAAAAAAAAAAAAAA96555550E542A96155101AFFFF953FFFFAE6A;
defparam sdpb_inst_14.INIT_RAM_0D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9566A561;
defparam sdpb_inst_14.INIT_RAM_0E = 256'h4516AAAAAAAAAAAAAAAAAAAAAAAAAAAA955550F546A961058C6AFFE44BFFFFEA;
defparam sdpb_inst_14.INIT_RAM_0F = 256'hEA6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5;
defparam sdpb_inst_14.INIT_RAM_10 = 256'hA9555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA655550250AA97D5151ABFE56FFFFF;
defparam sdpb_inst_14.INIT_RAM_11 = 256'hFFEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_12 = 256'hAAA9555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5554250AA9741206BFD13FFF;
defparam sdpb_inst_14.INIT_RAM_13 = 256'hFFFFEA6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_14 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95550E51AA578486AA54FF;
defparam sdpb_inst_14.INIT_RAM_15 = 256'hFFFFFFAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_16 = 256'hAAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAA6AAAAAAAAAAAAA5550E51AA415319552;
defparam sdpb_inst_14.INIT_RAM_17 = 256'h2FEFFFFFAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_18 = 256'hAAAAAAAAAAAA9AAAAAAAA66AAAA9AAAAAAAAAAAAAAAAAAAAA5550E52AA559854;
defparam sdpb_inst_14.INIT_RAM_19 = 256'h27FFFFFFFEA96AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA6AAAAAA;
defparam sdpb_inst_14.INIT_RAM_1A = 256'h69AAA6A5A695AAAAA9A9A9AAAAAAAA9AAAAAAAAAAAAAAAAAAAAA5550D52A75A7;
defparam sdpb_inst_14.INIT_RAM_1B = 256'h5AFFFFFEFFFFA5AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AA565A9;
defparam sdpb_inst_14.INIT_RAM_1C = 256'h6565665555555AAA5A665A5AAAAA5A959AAAAAAAA6AAAAAAAAAAAAA5540E56A5;
defparam sdpb_inst_14.INIT_RAM_1D = 256'h295A0FFFFEFFEAD5AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA96669;
defparam sdpb_inst_14.INIT_RAM_1E = 256'h5955555555555556A55A6656656A56A556699996AAAAAAAAAAAAAAAAAA5543E4;
defparam sdpb_inst_14.INIT_RAM_1F = 256'h3E40656FFFFF3FFEA5AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95A555;
defparam sdpb_inst_14.INIT_RAM_20 = 256'h556555555555555559555555555555555555555565599AAAAAAAAAAAAAAA9554;
defparam sdpb_inst_14.INIT_RAM_21 = 256'h5503E58456FFFB0BEB56AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555;
defparam sdpb_inst_14.INIT_RAM_22 = 256'h555555555555555555555555555555555555555555555559AAAAAAAAAAAAAAA9;
defparam sdpb_inst_14.INIT_RAM_23 = 256'hAA95503E1D35AFFBF2AD56AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA955;
defparam sdpb_inst_14.INIT_RAM_24 = 256'h5555555555555555555555555555555555555555555555656566AAAAAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_25 = 256'hAAAAA95503E0A2BA1FFCAB5AAAAAAAAAAAAAAAAAA6AAAAA6A669A9AA9AA6A955;
defparam sdpb_inst_14.INIT_RAM_26 = 256'h55555555555555555555555555555555555555555555555555555AAAAAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_27 = 256'hAAAAAAAA55503E562FA5FDAD56AAAAAAAAAAAAAAA9955A6A55655696A595AAA5;
defparam sdpb_inst_14.INIT_RAM_28 = 256'h95555555555555555555555555555555555555555555555555555556AAAAAAAA;
defparam sdpb_inst_14.INIT_RAM_29 = 256'hAAAAAAAAAAA55543E5DAF3F8B56AAAAAAAAAAAAAAAA955555555555555555555;
defparam sdpb_inst_14.INIT_RAM_2A = 256'h55555555555555555555555555555555555555555555555555555555556AAAAA;
defparam sdpb_inst_14.INIT_RAM_2B = 256'hAAAAAAAAAAAAAA55543FABFFFA15AAAAAAAAAAAAAAAAA6555555555555555555;
defparam sdpb_inst_14.INIT_RAM_2C = 256'h555555555555555555555555555555555555555555555555555555555555556A;
defparam sdpb_inst_14.INIT_RAM_2D = 256'h5AAAAAAAAAAAAAAAA9555003FC05556AAAAAAAAAAAAAAA655555555555555555;
defparam sdpb_inst_14.INIT_RAM_2E = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sdpb_inst_14.INIT_RAM_2F = 256'h555A6AAAAAAAAAAAAAAA955554055556AAAAAAAAAAAAAAA99955555555555555;
defparam sdpb_inst_14.INIT_RAM_30 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sdpb_inst_14.INIT_RAM_31 = 256'h5555555AAAAAAAAAAAAAAAA9555555555AAAAAAAAAAAAAAAA555555555555555;
defparam sdpb_inst_14.INIT_RAM_32 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam sdpb_inst_14.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000155555555;

SDPB sdpb_inst_15 (
    .DO({sdpb_inst_15_dout_w[30:0],sdpb_inst_15_dout[6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[6]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_15.READ_MODE = 1'b1;
defparam sdpb_inst_15.BIT_WIDTH_0 = 1;
defparam sdpb_inst_15.BIT_WIDTH_1 = 1;
defparam sdpb_inst_15.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_15.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_15.RESET_MODE = "SYNC";
defparam sdpb_inst_15.INIT_RAM_00 = 256'h000000000000000000DFEFFFFFFFE40000000000008002020000000000000002;
defparam sdpb_inst_15.INIT_RAM_01 = 256'h0000000000000000001DFFF3FFFFF650000000000000901C5000000000000000;
defparam sdpb_inst_15.INIT_RAM_02 = 256'h00000000000000000002FFFDEFFFFFFD408000008479F3FC3A20000000000000;
defparam sdpb_inst_15.INIT_RAM_03 = 256'h00000000000000000005F7FF3FFFFFFF9C8100057DFD7FFB79E3048000000000;
defparam sdpb_inst_15.INIT_RAM_04 = 256'h000000000000000000007BFFCFFFFFFFBFEF0FA36FFFFFFFEE3BBF8000000000;
defparam sdpb_inst_15.INIT_RAM_05 = 256'h0000000000000000000001FFFDFFE0FFFEFF88D4FF4DFFFFFEEABFE000000000;
defparam sdpb_inst_15.INIT_RAM_06 = 256'h0000000000000000000010FFFF07F877FFFFB8C5E79BFFFFFFFFC7F910000000;
defparam sdpb_inst_15.INIT_RAM_07 = 256'h000000000000000000000007DF9E1F1FCFFBF24065F9FFFFFFFF6F91A5800000;
defparam sdpb_inst_15.INIT_RAM_08 = 256'h0000000000000000000000017FFBF843FF7FE3E805AFFFFFFFFFFEFF88800000;
defparam sdpb_inst_15.INIT_RAM_09 = 256'h00000000000000000000000003FCFFE0FFF801160084F9FFBFFF7FF7FF420000;
defparam sdpb_inst_15.INIT_RAM_0A = 256'h00000000000000000000000001BFDFFE67FE380048804B7FABF4FFFFBE840904;
defparam sdpb_inst_15.INIT_RAM_0B = 256'h0000000000000000000000000017D8FF861FC7E00000007FFFFFDCAFFFD01250;
defparam sdpb_inst_15.INIT_RAM_0C = 256'h8E01006000000000000000000000DDC3F0F871FF8000020FFFFFFF4AFFFF9112;
defparam sdpb_inst_15.INIT_RAM_0D = 256'h1000000000000000000000000000A3BF0C3FE03FFC000001FFFF83EFFF7EFB90;
defparam sdpb_inst_15.INIT_RAM_0E = 256'h9020000000000000000000000000000FFC0FFF83FF8000001FEFC3E3D717FFB0;
defparam sdpb_inst_15.INIT_RAM_0F = 256'h582400C0000000000000000000000053FFE0FFF00FE2000005FFF1D50FFF4FDC;
defparam sdpb_inst_15.INIT_RAM_10 = 256'hFF31E10D6000040000000000000000003FFC03FC3C3C000000FFFCFBBCFFFEFF;
defparam sdpb_inst_15.INIT_RAM_11 = 256'hFFF8800004000200000000000000000000FF0E0F8FF00000000BBFDFD1C5FFFF;
defparam sdpb_inst_15.INIT_RAM_12 = 256'hFFFFF5800810100204000000000000000043E3F821FFC0000000DFF1E1E00FFF;
defparam sdpb_inst_15.INIT_RAM_13 = 256'hFFFFFFFC4024006800000000000000000010087FE27FFC0000000FF90E70007F;
defparam sdpb_inst_15.INIT_RAM_14 = 256'h1FFE77FE8100200800000000000000000000041FFF33FF880000027BD0740023;
defparam sdpb_inst_15.INIT_RAM_15 = 256'h71FFE0FFFFC09201000020000000000000000011FFE00FE00000000FFF038006;
defparam sdpb_inst_15.INIT_RAM_16 = 256'h7B87FCFB73E84001C3600800000000000000002007F8783C080000007FF81000;
defparam sdpb_inst_15.INIT_RAM_17 = 256'h7EF47FFFFF204000088200000000000000000000081F1FE0108A000001FE8083;
defparam sdpb_inst_15.INIT_RAM_18 = 256'h2373E1FFFFFFF804385C7008000000000000000000A043FF800A0000008BF004;
defparam sdpb_inst_15.INIT_RAM_19 = 256'h005ED70FFFFFE3AC10991AA80000000000000000000200FFFC00800000010000;
defparam sdpb_inst_15.INIT_RAM_1A = 256'h0002F3CCBFFFFEBE00821C8A0400000000000000000D4007FF08080000000000;
defparam sdpb_inst_15.INIT_RAM_1B = 256'h00801EF7E3FFFFFF040213C55010000000000000000091041FE0810000000000;
defparam sdpb_inst_15.INIT_RAM_1C = 256'hC00000FF9F1FFFFDE0080018890080000000000000000010007C880000000000;
defparam sdpb_inst_15.INIT_RAM_1D = 256'h00000007E6B87FFFFF000400E704000000000000000000020001008A00000001;
defparam sdpb_inst_15.INIT_RAM_1E = 256'h0407C0003FAF43FFFFDC44000C82020000000000000000042C00040800600000;
defparam sdpb_inst_15.INIT_RAM_1F = 256'h0002038001F73E0FDFFD860007F4E90000000000000000002002000000000000;
defparam sdpb_inst_15.INIT_RAM_20 = 256'h00108003020FED705FEFF008443B46000000000000002C000090000000020000;
defparam sdpb_inst_15.INIT_RAM_21 = 256'h000210000C007F5E8197FE100042D2C900000000000004000013424140004000;
defparam sdpb_inst_15.INIT_RAM_22 = 256'h00000200002003EE7C037FF03000055800000000000040422000401010040200;
defparam sdpb_inst_15.INIT_RAM_23 = 256'h000000200001000FDAF00C2B00104184904000000000000022001120000A4000;
defparam sdpb_inst_15.INIT_RAM_24 = 256'h0800004400000C007FBC0042C00000103E800000000020801400000004200440;
defparam sdpb_inst_15.INIT_RAM_25 = 256'h840000000000004003DF0000029008535BEC0000000000202000000020841004;
defparam sdpb_inst_15.INIT_RAM_26 = 256'h1040000044000002001FE0C000000A00425A0000000000010000200044181204;
defparam sdpb_inst_15.INIT_RAM_27 = 256'h03000000040000002000F0200000050829B38200000000000000008001102080;
defparam sdpb_inst_15.INIT_RAM_28 = 256'h00B100000040000002200C00000080020010808000000000000000000007000A;
defparam sdpb_inst_15.INIT_RAM_29 = 256'hA0412000000210000000006000000400801B1330000000000000000000001048;
defparam sdpb_inst_15.INIT_RAM_2A = 256'h0088000000002000000020020000000000237E6C600000000000000000000001;
defparam sdpb_inst_15.INIT_RAM_2B = 256'h0200020000000100000004003000000000400288E00000000000000000C00000;
defparam sdpb_inst_15.INIT_RAM_2C = 256'h0020002000000018400010000200000000000C33BB4C00000000000100000000;
defparam sdpb_inst_15.INIT_RAM_2D = 256'h00000204000000008000000000300000000004541FED40000000000000000000;
defparam sdpb_inst_15.INIT_RAM_2E = 256'h00000200800000000400000000030000000000000BC390000000000000000100;
defparam sdpb_inst_15.INIT_RAM_2F = 256'h00000000800000000060000000003000000000084137AE000000000000000000;
defparam sdpb_inst_15.INIT_RAM_30 = 256'h0000000004000000000200001800018000000000204F17500000000000000000;
defparam sdpb_inst_15.INIT_RAM_31 = 256'h0080000000000000000010000600001C0000000000117D288000000000000000;
defparam sdpb_inst_15.INIT_RAM_32 = 256'h0018000000000000000000E011000000C000000000061147A000000000000200;
defparam sdpb_inst_15.INIT_RAM_33 = 256'h00018000000000000000000131C00000060000020008021FFC20000000000000;
defparam sdpb_inst_15.INIT_RAM_34 = 256'h1000DC000000000000000000001000000038000020000CECFF80000000000001;
defparam sdpb_inst_15.INIT_RAM_35 = 256'h00007F800000000000000000000000000001C0001A00000D2BF4000000000000;
defparam sdpb_inst_15.INIT_RAM_36 = 256'h0000FFF80000000000000000000000000800060007F00008990FC80000000000;
defparam sdpb_inst_15.INIT_RAM_37 = 256'h000000C70000000000000000000000000200003E01FE80020239440000000000;
defparam sdpb_inst_15.INIT_RAM_38 = 256'h00000024E00000000000000000000000000000003C1F9C000091F03800000000;
defparam sdpb_inst_15.INIT_RAM_39 = 256'h000000013C0000000000000000000000000100000027E7A00019493600000000;
defparam sdpb_inst_15.INIT_RAM_3A = 256'h0000000004000000000000000000000000000280000175E70080B15FE0000000;
defparam sdpb_inst_15.INIT_RAM_3B = 256'h000000000000000000000000000000000000000400000BF9F817024479400000;
defparam sdpb_inst_15.INIT_RAM_3C = 256'h00000000000000000000000000000000000000000000007DFBC2B034C7900000;
defparam sdpb_inst_15.INIT_RAM_3D = 256'h0000000000000004000000000000000000001CC000000003FA76101000F41000;
defparam sdpb_inst_15.INIT_RAM_3E = 256'h0000000000000000600000000000000000003C00000000001EFAF000408DD800;
defparam sdpb_inst_15.INIT_RAM_3F = 256'h000000000000000004C00000000000000000FC000000000000FE9D848498C400;

SDPB sdpb_inst_16 (
    .DO({sdpb_inst_16_dout_w[30:0],sdpb_inst_16_dout[6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[6]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_16.READ_MODE = 1'b1;
defparam sdpb_inst_16.BIT_WIDTH_0 = 1;
defparam sdpb_inst_16.BIT_WIDTH_1 = 1;
defparam sdpb_inst_16.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_16.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_16.RESET_MODE = "SYNC";
defparam sdpb_inst_16.INIT_RAM_00 = 256'h000000000000000000D9000010000000001FF000000000000007BEBC08001C88;
defparam sdpb_inst_16.INIT_RAM_01 = 256'hD000000000000000003B100002001000003C00000000000000003FA7E0002398;
defparam sdpb_inst_16.INIT_RAM_02 = 256'h26000000000000000005430000000080003C000000000000000001EFBE000002;
defparam sdpb_inst_16.INIT_RAM_03 = 256'h24400000000000000000252000000000001E000000000000C000000FCB300010;
defparam sdpb_inst_16.INIT_RAM_04 = 256'h04280000000000000000008400000000000F000000100000008000007BCF8000;
defparam sdpb_inst_16.INIT_RAM_05 = 256'h0108800000000000000000408000000008030000008700000700000003F2DC00;
defparam sdpb_inst_16.INIT_RAM_06 = 256'h000058000000000000000010300000000000C0000018000000000000001EF3E0;
defparam sdpb_inst_16.INIT_RAM_07 = 256'hF80020000000000000000000060000020020600000580000000000200000FCB7;
defparam sdpb_inst_16.INIT_RAM_08 = 256'h2DC00028000000000000000000C00000000408000004000000000000600007FC;
defparam sdpb_inst_16.INIT_RAM_09 = 256'hFF3F000C0000000000000000001800000100830000020000000000000020003F;
defparam sdpb_inst_16.INIT_RAM_0A = 256'h0FCB7800000000000000000000090000000020C0000080000000000000048001;
defparam sdpb_inst_16.INIT_RAM_0B = 256'h007FCFC000000000000000000010300000004810000140000000000000008000;
defparam sdpb_inst_16.INIT_RAM_0C = 256'h0003F2CE00080000000000000002060000000006000010000000000000000080;
defparam sdpb_inst_16.INIT_RAM_0D = 256'h00001FF3F000800000000000000000C000000000C00000000000000000000000;
defparam sdpb_inst_16.INIT_RAM_0E = 256'h000000FCB3800000000000000000000800000000080000000000000000000000;
defparam sdpb_inst_16.INIT_RAM_0F = 256'h00000007FCF40030000000000000000180000000010000000000000000000000;
defparam sdpb_inst_16.INIT_RAM_10 = 256'h000000003F2CE0000000000000000010B0000000002000100000000000000000;
defparam sdpb_inst_16.INIT_RAM_11 = 256'h0000000001FF3D00000000000000000222000000000400000000000000000000;
defparam sdpb_inst_16.INIT_RAM_12 = 256'h000000000007CB380000000000000000006000000000C0000000000000000000;
defparam sdpb_inst_16.INIT_RAM_13 = 256'h0000000000007BCF4000000000000000000C0000000018000000000000000000;
defparam sdpb_inst_16.INIT_RAM_14 = 256'h00000000000001F2CE0000000000000000058000000001000000000000000000;
defparam sdpb_inst_16.INIT_RAM_15 = 256'h0000000000000006F3D000000000000000041800000000200000000000000000;
defparam sdpb_inst_16.INIT_RAM_16 = 256'h00000000000000007C9B80000000000000020300000000040004000000000000;
defparam sdpb_inst_16.INIT_RAM_17 = 256'h000000000000000003BEFC00000000000000416000000000C001000000000000;
defparam sdpb_inst_16.INIT_RAM_18 = 256'h0000000000000000001FA6E00000000000000024000000000800000000000000;
defparam sdpb_inst_16.INIT_RAM_19 = 256'h000000000000000000006B8F800000000001F000C00000000100000000000000;
defparam sdpb_inst_16.INIT_RAM_1A = 256'h0000000000000000000007EDAC0000000000FFE0180000000030002000000000;
defparam sdpb_inst_16.INIT_RAM_1B = 256'h00000000000000000000001A7DE0000000001FF80B8000000002000000000000;
defparam sdpb_inst_16.INIT_RAM_1C = 256'h000000000000000000000000FB7B0000000007FF90B000000000200000000000;
defparam sdpb_inst_16.INIT_RAM_1D = 256'h0000000000000000000000000E9F78000000007FF03F00000000040018000000;
defparam sdpb_inst_16.INIT_RAM_1E = 256'h000000000000000000000000007FCEC00000000FFE07F800000000C000000000;
defparam sdpb_inst_16.INIT_RAM_1F = 256'h0000000000040000000000000003E7DE00000001FF003FE00000000800000000;
defparam sdpb_inst_16.INIT_RAM_20 = 256'h00000000000004000000000000001FF3900000001FC007FC0000000180000000;
defparam sdpb_inst_16.INIT_RAM_21 = 256'h0000000000178004000000000000007D2380000001F8007FF000000010000000;
defparam sdpb_inst_16.INIT_RAM_22 = 256'h000000000006FF0000000000000000077CFC0000003F8003FE80000003000000;
defparam sdpb_inst_16.INIT_RAM_23 = 256'h0000000000019FFC00000000000000000F2FC0000003F8013FC80000002000C0;
defparam sdpb_inst_16.INIT_RAM_24 = 256'h0000000000002FFFF00000000000000000CBFC000000670007FD800000020000;
defparam sdpb_inst_16.INIT_RAM_25 = 256'h00000000000005FFFFC00000000000000003FFC000001B7900FF900000006000;
defparam sdpb_inst_16.INIT_RAM_26 = 256'h01000000000000BFFFFE00000000000000003FFC000006FF851FFB0000000200;
defparam sdpb_inst_16.INIT_RAM_27 = 256'h0000000000000017FFFFF80000000000000002FF80000187FE03FF2000000040;
defparam sdpb_inst_16.INIT_RAM_28 = 256'h4000000000000002FFFFFFE0000000000000000FF0000063FFFFFFC400000004;
defparam sdpb_inst_16.INIT_RAM_29 = 256'h0C000000000000007FFE3FFB80000000000000000000000C7BFFFFF980000000;
defparam sdpb_inst_16.INIT_RAM_2A = 256'h008000000000000005FFC0BF9E0000000000000000000003DC7FFFFF30000000;
defparam sdpb_inst_16.INIT_RAM_2B = 256'h000800000000000000BFF807F870000000000000000000007F83FFFFE7000000;
defparam sdpb_inst_16.INIT_RAM_2C = 256'h00008003000000000017FF001FC3C00000000000000000000FF17FEFFCE00000;
defparam sdpb_inst_16.INIT_RAM_2D = 256'h000018000000000000037FF0007F0300000000000000000001FC03FEFFDC0000;
defparam sdpb_inst_16.INIT_RAM_2E = 256'h0000010000000000000027FE0000FC0C0000000000000000003F802FC1FDC000;
defparam sdpb_inst_16.INIT_RAM_2F = 256'h000000100000000000000279400003F060000000000000000000E3009803D800;
defparam sdpb_inst_16.INIT_RAM_30 = 256'h0000000100060000000000C7FC00003F89800000000000000000407781003D80;
defparam sdpb_inst_16.INIT_RAM_31 = 256'h800000001000000000000004FF800003FEE60000000000000000001FFC0003D8;
defparam sdpb_inst_16.INIT_RAM_32 = 256'hD800000001000000000000018FFE00007FFFB0000000000000000000FFF8003D;
defparam sdpb_inst_16.INIT_RAM_33 = 256'h0D800000002000000000000019F7F8000FFFFCC00000000000000008008FFC01;
defparam sdpb_inst_16.INIT_RAM_34 = 256'h00980000000000000000000001FEB3A0003BFFF3000000000000000080000380;
defparam sdpb_inst_16.INIT_RAM_35 = 256'h000180000000200000000000001FE68CC00287FF4C0000000000000000000000;
defparam sdpb_inst_16.INIT_RAM_36 = 256'h0000300000000200000000000001FFFF3302100FF60000000000000000400000;
defparam sdpb_inst_16.INIT_RAM_37 = 256'h00008300000000600000000000001FFFFE4442000F0C40000000000000000000;
defparam sdpb_inst_16.INIT_RAM_38 = 256'h000024600000000400000000000000FFFFFD100000E03B000000000000002000;
defparam sdpb_inst_16.INIT_RAM_39 = 256'h1800030C0000000040020000000000073FDFF7640006007C0000000000000100;
defparam sdpb_inst_16.INIT_RAM_3A = 256'h217401C0C0000000040000000000000072FFFE798000E001F000000000000008;
defparam sdpb_inst_16.INIT_RAM_3B = 256'h0082BCE038000000014000000000000003C3FF01E0000C000F80000000000000;
defparam sdpb_inst_16.INIT_RAM_3C = 256'h000300C0060000000000002000000000001E0FE00780008000FE000000000000;
defparam sdpb_inst_16.INIT_RAM_3D = 256'h00000E0001C0000000002002000000000000717F801E00380007F00000000000;
defparam sdpb_inst_16.INIT_RAM_3E = 256'h0000001B887000000000060040000000000003C3FC00B80100007F8000000000;
defparam sdpb_inst_16.INIT_RAM_3F = 256'h000000003FF8000000000240040000000000000FDFF800C0100007E800000000;

SDPB sdpb_inst_17 (
    .DO({sdpb_inst_17_dout_w[30:0],sdpb_inst_17_dout[7]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_17.READ_MODE = 1'b1;
defparam sdpb_inst_17.BIT_WIDTH_0 = 1;
defparam sdpb_inst_17.BIT_WIDTH_1 = 1;
defparam sdpb_inst_17.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_17.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_17.RESET_MODE = "SYNC";
defparam sdpb_inst_17.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_17.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8078FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE1E0E03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFC07BC00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF001F0007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0019801C7FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0079E0381FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3C0F078E007FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0F3C01FC003FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003F0007C007FFFFFFFFFFC1FFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC001F000FF01CFFFFFFFFFE20FFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC003FC03C3C38FFFFFFFFF0043FFFFFF;
defparam sdpb_inst_17.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00F1F0700FF0FFFFFFFFE02E3FFFFF;
defparam sdpb_inst_17.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBC1C07DE003C0FFFFFFFFE1E007FFF;
defparam sdpb_inst_17.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F7801F8003C0FFFFFFFFF18003FF;
defparam sdpb_inst_17.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3E000CC00740FFFFFFFFF80001F;
defparam sdpb_inst_17.INIT_RAM_15 = 256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0E001FF01CC1FFFFFFFFFC0001;
defparam sdpb_inst_17.INIT_RAM_16 = 256'h007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0F80787C3843FFFFFFFFFE000;
defparam sdpb_inst_17.INIT_RAM_17 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE05E0E01FE044FFFFFFFFFF00;
defparam sdpb_inst_17.INIT_RAM_18 = 256'hC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF047BC007C058FFFFFFFFFF8;
defparam sdpb_inst_17.INIT_RAM_19 = 256'hFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC41F0003C070FFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_1A = 256'hFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2207800E4060FFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_1B = 256'h427FE0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0E03E01C40C0FFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_1C = 256'h0003FF0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF860378304340FFFFFFC;
defparam sdpb_inst_17.INIT_RAM_1D = 256'hC00007F80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81831EE04441FFFFFE;
defparam sdpb_inst_17.INIT_RAM_1E = 256'hF8000007C0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF812307807840FFFFF;
defparam sdpb_inst_17.INIT_RAM_1F = 256'hFF01FC007E0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC19901807048FFFF;
defparam sdpb_inst_17.INIT_RAM_20 = 256'hFFE07FFC01F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFF0878180E050FFF;
defparam sdpb_inst_17.INIT_RAM_21 = 256'hFFFC0FFFF00F80007FFFFFFFFFFFFFFFFFFFFFFFFFF8F83FFFEC818081E020FF;
defparam sdpb_inst_17.INIT_RAM_22 = 256'hFFFFC1FFFFC0FC0003FFFFFFFFFFFFFFFFFFFFFFFFFF0781C3FE3C0E0C320C0F;
defparam sdpb_inst_17.INIT_RAM_23 = 256'h3FFFFC1FFFFE03F0000FFFFFFFFFFFFFFFFFFFFFFFFFF07C1C1FE0C0B8C42161;
defparam sdpb_inst_17.INIT_RAM_24 = 256'h67FFFF83FFFFF03F8000003FFFFFFFFFFFFFFFFFFFFFC307E3C1FF0708CD8226;
defparam sdpb_inst_17.INIT_RAM_25 = 256'h03FFFFF83FFFFF83FC000000FFFFFFFFFFFFFFFFFFFFFC1E1F3E3FF05C43E068;
defparam sdpb_inst_17.INIT_RAM_26 = 256'h603FFFFF83FFFFFC1FE0000003FFFFFFFFFFFFFFFFFFFFC0F0F1C7FF82640C03;
defparam sdpb_inst_17.INIT_RAM_27 = 256'h0C07FFFFF83FFFFFC1FF0000001FFFFFFFFFFFFFFFFFFFFE0380007FFE21C040;
defparam sdpb_inst_17.INIT_RAM_28 = 256'h6100FFFFFF83FFFFFC1FF00000007FFFFFFFFFFFFFFFFFFFFC00000FFFF80604;
defparam sdpb_inst_17.INIT_RAM_29 = 256'h46221FFFFFFC0FFFFFC1FF80000003FFFFFFFFFFFFFFFFFFFFF00000FFFFE030;
defparam sdpb_inst_17.INIT_RAM_2A = 256'h336437FFFFFFC0FFFFF81FFC0000003FFFFFFFFFFFFFFFFFFFFF80000FFFFF82;
defparam sdpb_inst_17.INIT_RAM_2B = 256'hF90F81FFFFFFFE07FFFF03FFC0000001FFFFFFFFFFFFFFFFFFFFFE00003FFFFE;
defparam sdpb_inst_17.INIT_RAM_2C = 256'hFFD0301FFFFFFFE03FFFE07FFC0000001FFFFFFFFFFFFFFFFFFFFFFE0003FFFF;
defparam sdpb_inst_17.INIT_RAM_2D = 256'hFFFF8103FFFFFFFF03FFFC0FFFC0000001FFFFFFFFFFFFFFFFFFFFFFE0001FFF;
defparam sdpb_inst_17.INIT_RAM_2E = 256'hFFFFFC107FFFFFFFF81FFE01FFFC0000001FFFFFFFFFFFFFFFFFFFFFFC0000FF;
defparam sdpb_inst_17.INIT_RAM_2F = 256'h7FFFFFF11FFFFFFFFF81FF003FFFC0000001FFFFFFFFFFFFFFFFFFFFFFC0000F;
defparam sdpb_inst_17.INIT_RAM_30 = 256'h07FFFFFFDBFFFFFFFFFC010007FFFE0000001FFFFFFFFFFFFFFFFFFFFFFC0000;
defparam sdpb_inst_17.INIT_RAM_31 = 256'h007FFFFFFFFFFFFFFFFFE00001FFFFE0000001FFFFFFFFFFFFFFFFFFFFFFC000;
defparam sdpb_inst_17.INIT_RAM_32 = 256'h0007FFFFFFFFFFFFFFFFFF0000FFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_17.INIT_RAM_33 = 256'h00007FFFFFFFFFFFFFFFFFFE003FFFFFF8000001FFFFFFFFFFFFFFFFFFFFFFE0;
defparam sdpb_inst_17.INIT_RAM_34 = 256'hE00003FFFFFFFFFFFFFFFFFFFFEFFFFFFFC000001FFFFFFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_17.INIT_RAM_35 = 256'hFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000001FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_36 = 256'hFFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_37 = 256'hFFFFFF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_38 = 256'hFFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_39 = 256'hFFFFFFFE03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_3A = 256'hFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFF00007FFFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC07FFFFFFF80003FFFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFF8FFFFFFFFFFFFFFFFFFFFE03FFFFFFFFC0001FFFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFF01FFFFFFFFFFFFFFFFFFC3FFFFFFFFFFE0000FFFFFFFFFFF;
defparam sdpb_inst_17.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFFF03FFFFFFFFFFFF00007FFFFFFFFF;

SDPB sdpb_inst_18 (
    .DO({sdpb_inst_18_dout_w[30:0],sdpb_inst_18_dout[7]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[15],ada[14]}),
    .BLKSELB({gw_gnd,adb[15],adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_18.READ_MODE = 1'b1;
defparam sdpb_inst_18.BIT_WIDTH_0 = 1;
defparam sdpb_inst_18.BIT_WIDTH_1 = 1;
defparam sdpb_inst_18.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_18.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_18.RESET_MODE = "SYNC";
defparam sdpb_inst_18.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFE00FFFFE007FFFFFFE00FFFFFFFFFFFFFF80003FFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFC00FFFFC000FFFFFC3FFFFFFFFFFFFFFFFC0001FFFFFFF;
defparam sdpb_inst_18.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFF820FFFFC0007FFFC3FFFFFFFFFFFFFFFFFE0001FFFFFF;
defparam sdpb_inst_18.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFF801FFFFC0007FFE1FFFFFFFFFFFF07FFFFF0000FFFFF;
defparam sdpb_inst_18.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFF803FFFFC0007FF0FFFFFFE00000007FFFFF80007FFF;
defparam sdpb_inst_18.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFF007FFFFC0007FCFFFFFF00FFFFF8FFFFFFFC0003FF;
defparam sdpb_inst_18.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFE00FFFFFC000FF3FFFFF07FFFFFFFFFFFFFFE0001F;
defparam sdpb_inst_18.INIT_RAM_07 = 256'h07FFFFFFFFFFFFFFFFFFFFFE01FFFFFC001F9FFFFF87FFFFFFFFFFFFFFFF0000;
defparam sdpb_inst_18.INIT_RAM_08 = 256'h003FFFFFFFFFFFFFFFFFFFFFC03FFFFFE003F7FFFFE3FFFFFFFFFFFFFFFFF800;
defparam sdpb_inst_18.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFFFFFFFF807FFFFFE007CFFFFF1FFFFFFFFFFFFFFFFFFC0;
defparam sdpb_inst_18.INIT_RAM_0A = 256'hF00007FFFFFFFFFFFFFFFFFFFF00FFFFFFF01F3FFFFC7FFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_18.INIT_RAM_0B = 256'hFF80003FFFFFFFFFFFFFFFFFFFE00FFFFFFF87EFFFFE3FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_0C = 256'hFFFC0001FFFFFFFFFFFFFFFFFFFC01FFFFFFFFF9FFFF8FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_0D = 256'hFFFFE0000FFFFFFFFFFFFFFFFFFFC03FFFFFFFFF3FFFE7FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_0E = 256'hFFFFFF00007FFFFFFFFFFFFFFFFFF807FFFFFFFFF7FFF9FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_0F = 256'hFFFFFFF80003FFFFFFFFFFFFFFFFFF007FFFFFFFFEFFFE7FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_10 = 256'hFFFFFFFFC0001FFFFFFFFFFFFFFFFFE00FFFFFFFFFDFFFCFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_11 = 256'hFFFFFFFFFE0000FFFFFFFFFFFFFFFFFC01FFFFFFFFFBFFFBFFFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_12 = 256'hFFFFFFFFFFF80007FFFFFFFFFFFFFFFFC01FFFFFFFFF3FFF7FFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_13 = 256'hFFFFFFFFFFFF80003FFFFFFFFFFFFFFFF803FFFFFFFFE7FFEFFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_14 = 256'hFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFF007FFFFFFFFEFFFDFFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFE007FFFFFFFFDFFFBFFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFC00FFFFFFFFFBFFF3FFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFF801FFFFFFFFF3FFE7FFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFF803FFFFFFFFF7FFEFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFF00007FFFFFFFFFFE0F003FFFFFFFFEFFFDFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFF000007FFFFFFFFCFFF9FFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFC0001FFFFFFFFFE000007FFFFFFFFDFFFBFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFE0000FFFFFFFFF800000FFFFFFFFF9FFF7FFFFFFF;
defparam sdpb_inst_18.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF00007FFFFFFFF800000FFFFFFFFFBFFE7FFFFFF;
defparam sdpb_inst_18.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFF0000007FFFFFFFF3FFEFFFFFF;
defparam sdpb_inst_18.INIT_RAM_1F = 256'hFFFFFFFFFFFBFFFFFFFFFFFFFFFC0001FFFFFFFE0000001FFFFFFFF7FFDFFFFF;
defparam sdpb_inst_18.INIT_RAM_20 = 256'hFFFFFFFFFFFFFBFFFFFFFFFFFFFFE0000FFFFFFFE0000001FFFFFFFE7FFDFFFF;
defparam sdpb_inst_18.INIT_RAM_21 = 256'hFFFFFFFFFFE07FFBFFFFFFFFFFFFFF00007FFFFFFE0000000FFFFFFFEFFFBFFF;
defparam sdpb_inst_18.INIT_RAM_22 = 256'hFFFFFFFFFFF800FFFFFFFFFFFFFFFFF80003FFFFFFC00000007FFFFFFCFFFBFF;
defparam sdpb_inst_18.INIT_RAM_23 = 256'hFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFC0003FFFFFFC00000007FFFFFFDFFF3F;
defparam sdpb_inst_18.INIT_RAM_24 = 256'h7FFFFFFFFFFFC0000FFFFFFFFFFFFFFFFE0003FFFFFF800000007FFFFFFDFFF7;
defparam sdpb_inst_18.INIT_RAM_25 = 256'hF7FFFFFFFFFFF800003FFFFFFFFFFFFFFFF0003FFFFFE40000000FFFFFFF9FFF;
defparam sdpb_inst_18.INIT_RAM_26 = 256'hFEFFFFFFFFFFFF000001FFFFFFFFFFFFFFFF8003FFFFF900000000FFFFFFF9FF;
defparam sdpb_inst_18.INIT_RAM_27 = 256'hFFEFFFFFFFFFFFE0000007FFFFFFFFFFFFFFFC007FFFFE780000001FFFFFFFBF;
defparam sdpb_inst_18.INIT_RAM_28 = 256'hBFFEFFFFFFFFFFFC0000001FFFFFFFFFFFFFFFF00FFFFF9C00000003FFFFFFFB;
defparam sdpb_inst_18.INIT_RAM_29 = 256'hF3FFEFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFF3840000007FFFFFFF;
defparam sdpb_inst_18.INIT_RAM_2A = 256'hFF7FFEFFFFFFFFFFF800004001FFFFFFFFFFFFFFFFFFFFFC200000000FFFFFFF;
defparam sdpb_inst_18.INIT_RAM_2B = 256'hFFF7FFEFFFFFFFFFFF000000000FFFFFFFFFFFFFFFFFFFFF8000000000FFFFFF;
defparam sdpb_inst_18.INIT_RAM_2C = 256'hFFFF7FFCFFFFFFFFFFE0000000003FFFFFFFFFFFFFFFFFFFF0000000001FFFFF;
defparam sdpb_inst_18.INIT_RAM_2D = 256'hFFFFE7FFDFFFFFFFFFFC0000000000FFFFFFFFFFFFFFFFFFFE0000000003FFFF;
defparam sdpb_inst_18.INIT_RAM_2E = 256'hFFFFFEFFFDFFFFFFFFFFC00000000003FFFFFFFFFFFFFFFFFFC0000000003FFF;
defparam sdpb_inst_18.INIT_RAM_2F = 256'hFFFFFFEFFFDFFFFFFFFFF806800000001FFFFFFFFFFFFFFFFFFC0000000007FF;
defparam sdpb_inst_18.INIT_RAM_30 = 256'hFFFFFFFEFFF9FFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFF80000000007F;
defparam sdpb_inst_18.INIT_RAM_31 = 256'h7FFFFFFFEFFFBFFFFFFFFFF0000000000001FFFFFFFFFFFFFFFFF80000000007;
defparam sdpb_inst_18.INIT_RAM_32 = 256'h07FFFFFFFEFFFBFFFFFFFFFE0000000000000FFFFFFFFFFFFFFFFF8000000000;
defparam sdpb_inst_18.INIT_RAM_33 = 256'h007FFFFFFFDFFFBFFFFFFFFFE00800000000003FFFFFFFFFFFFFFFF000000000;
defparam sdpb_inst_18.INIT_RAM_34 = 256'h0007FFFFFFFDFFF7FFFFFFFFFE014C4000C40000EFFFFFFFFFFFFFFF00000000;
defparam sdpb_inst_18.INIT_RAM_35 = 256'h00007FFFFFFFDFFF7FFFFFFFFFE01973001D780000FFFFFFFFFFFFFFF8000000;
defparam sdpb_inst_18.INIT_RAM_36 = 256'h00000FFFFFFFFDFFF7FFFFFFFFFE0000CC01EFF0000FFFFFFFFFFFFFFF800000;
defparam sdpb_inst_18.INIT_RAM_37 = 256'h000000FFFFFFFF9FFEFFFFFFFFFFE00001B83DFFF0003FFFFFFFFFFFFFFC0000;
defparam sdpb_inst_18.INIT_RAM_38 = 256'h0000001FFFFFFFFBFFEFFFFFFFFFFF000002E7FFFF0000FFFFFFFFFFFFFFC000;
defparam sdpb_inst_18.INIT_RAM_39 = 256'h00000003FFFFFFFFBFFCFFFFFFFFFFF80020089BFFF80003FFFFFFFFFFFFFE00;
defparam sdpb_inst_18.INIT_RAM_3A = 256'hC00000003FFFFFFFFBFFDFFFFFFFFFFF800000067FFF00000FFFFFFFFFFFFFF0;
defparam sdpb_inst_18.INIT_RAM_3B = 256'hFF00000007FFFFFFFE3FFDFFFFFFFFFFFC0000001FFFF000007FFFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_3C = 256'hFFFC000001FFFFFFFFE3FF9FFFFFFFFFFFE00000007FFF000001FFFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_3D = 256'hFFFFF000003FFFFFFFFE1FF9FFFFFFFFFFFF80000001FFC000000FFFFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_3E = 256'hFFFFFFE0000FFFFFFFFFE1FF3FFFFFFFFFFFFC00000007FE0000007FFFFFFFFF;
defparam sdpb_inst_18.INIT_RAM_3F = 256'hFFFFFFFFC007FFFFFFFFFC3FE3FFFFFFFFFFFFF00000003FE0000007FFFFFFFF;

SDPB sdpb_inst_19 (
    .DO({sdpb_inst_19_dout_w[29:0],sdpb_inst_19_dout[7:6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[15],ada[14],ada[13]}),
    .BLKSELB({adb[15],adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_19.READ_MODE = 1'b1;
defparam sdpb_inst_19.BIT_WIDTH_0 = 2;
defparam sdpb_inst_19.BIT_WIDTH_1 = 2;
defparam sdpb_inst_19.BLK_SEL_0 = 3'b100;
defparam sdpb_inst_19.BLK_SEL_1 = 3'b100;
defparam sdpb_inst_19.RESET_MODE = "SYNC";
defparam sdpb_inst_19.INIT_RAM_00 = 256'hAAAAAAAAAAAAAAAAA554555550000009AA940000000015545AAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_01 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA01AAAA81AAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_02 = 256'hAAAAAAAAAAAAAAAAAAAA55555555000001595000000000155456AAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_03 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA905AAAA81AAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_04 = 256'hAAAAAAAAAAAAAAAAAAAAAA95515555400000554000000000155455AAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_05 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA806AAAA41AAAAAAA;
defparam sdpb_inst_19.INIT_RAM_06 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAA9555555550000050000000000555565AAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_07 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5AAAAA41AAAAA;
defparam sdpb_inst_19.INIT_RAM_08 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555555590000100000000005555156AAAAA;
defparam sdpb_inst_19.INIT_RAM_09 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA06AAA;
defparam sdpb_inst_19.INIT_RAM_0A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA955455559000040000000015555516AAA;
defparam sdpb_inst_19.INIT_RAM_0B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA06A;
defparam sdpb_inst_19.INIT_RAM_0C = 256'h6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5555555800050000000015555556A;
defparam sdpb_inst_19.INIT_RAM_0D = 256'h6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA90;
defparam sdpb_inst_19.INIT_RAM_0E = 256'hA5AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555558001000000005555555;
defparam sdpb_inst_19.INIT_RAM_0F = 256'h556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_10 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95555554004000000055555;
defparam sdpb_inst_19.INIT_RAM_11 = 256'h55556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_12 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95555554010000001555;
defparam sdpb_inst_19.INIT_RAM_13 = 256'h555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_14 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555550040000055;
defparam sdpb_inst_19.INIT_RAM_15 = 256'h55555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_16 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555500100001;
defparam sdpb_inst_19.INIT_RAM_17 = 256'h1555555455AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_18 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555000400;
defparam sdpb_inst_19.INIT_RAM_19 = 256'h055555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_1A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55554544;
defparam sdpb_inst_19.INIT_RAM_1B = 256'h55555555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_1C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55555;
defparam sdpb_inst_19.INIT_RAM_1D = 256'h4555A5555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_1E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA955;
defparam sdpb_inst_19.INIT_RAM_1F = 256'h95544555555555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_20 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_21 = 256'hAAA9542055555495556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_22 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_23 = 256'hAAAAAA95555555415555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_24 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_25 = 256'hAAAAAAAAA9540065155555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_26 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_27 = 256'hAAAAAAAAAAAA955456915556AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_28 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_29 = 256'hAAAAAAAAAAAAAAA9551559055AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_2A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_2B = 256'hAAAAAAAAAAAAAAAAAA95555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_2C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_2D = 256'hAAAAAAAAAAAAAAAAAAAAAAA956AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_2E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_2F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_30 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_31 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_32 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_19.INIT_RAM_33 = 256'h00000000000000000000000000000000000000000000000000000002AAAAAAAA;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[15]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clkb),
  .CE(oce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clkb),
  .CE(oce)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_5 (
  .O(dout[0]),
  .I0(mux_o_3),
  .I1(sdpb_inst_4_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(sdpb_inst_2_dout[1]),
  .I1(sdpb_inst_3_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_11 (
  .O(dout[1]),
  .I0(mux_o_9),
  .I1(sdpb_inst_4_dout[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(sdpb_inst_5_dout[2]),
  .I1(sdpb_inst_6_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_17 (
  .O(dout[2]),
  .I0(mux_o_15),
  .I1(sdpb_inst_9_dout[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(sdpb_inst_7_dout[3]),
  .I1(sdpb_inst_8_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_23 (
  .O(dout[3]),
  .I0(mux_o_21),
  .I1(sdpb_inst_9_dout[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(sdpb_inst_10_dout[4]),
  .I1(sdpb_inst_11_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_29 (
  .O(dout[4]),
  .I0(mux_o_27),
  .I1(sdpb_inst_14_dout[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(sdpb_inst_12_dout[5]),
  .I1(sdpb_inst_13_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_35 (
  .O(dout[5]),
  .I0(mux_o_33),
  .I1(sdpb_inst_14_dout[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(sdpb_inst_15_dout[6]),
  .I1(sdpb_inst_16_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_41 (
  .O(dout[6]),
  .I0(mux_o_39),
  .I1(sdpb_inst_19_dout[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(sdpb_inst_17_dout[7]),
  .I1(sdpb_inst_18_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_47 (
  .O(dout[7]),
  .I0(mux_o_45),
  .I1(sdpb_inst_19_dout[7]),
  .S0(dff_q_1)
);
endmodule //Gowin_SDPB3
