//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Tue Aug 08 22:22:39 2023

module Gowin_SDPB4 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb); //488x302+1

output [0:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [17:0] ada;
input [0:0] din;
input [17:0] adb;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [0:0] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [0:0] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [0:0] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [0:0] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [0:0] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [0:0] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [0:0] sdpb_inst_7_dout;
wire [30:0] sdpb_inst_8_dout_w;
wire [0:0] sdpb_inst_8_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_5;
wire mux_o_6;
wire mux_o_8;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ada[14]),
  .I1(ada[15]),
  .I2(ada[16]),
  .I3(ada[17])
);
defparam lut_inst_8.INIT = 16'h0100;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_9.INIT = 16'h0001;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_10.INIT = 16'h0002;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_11.INIT = 16'h0004;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_12.INIT = 16'h0008;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_13.INIT = 16'h0010;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_14.INIT = 16'h0020;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_15.INIT = 16'h0040;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_16.INIT = 16'h0080;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(adb[14]),
  .I1(adb[15]),
  .I2(adb[16]),
  .I3(adb[17])
);
defparam lut_inst_17.INIT = 16'h0100;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_9}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00001FFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000007;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hFFFFFE000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFF0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FF;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam sdpb_inst_0.INIT_RAM_22 = 256'hFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_24 = 256'hFFFFFFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFE0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000007FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000003FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000003FFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000001FFFFF;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_0.INIT_RAM_37 = 256'hFFFFFE0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_1}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_10}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000001FFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000001FFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000FF;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000;
defparam sdpb_inst_1.INIT_RAM_0A = 256'hFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0C = 256'hFFFFFFFFC00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000001FFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000001FFFFF;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_1.INIT_RAM_1F = 256'hFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_21 = 256'hFFFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000003FFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000001FF;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam sdpb_inst_1.INIT_RAM_32 = 256'hFFC0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_34 = 256'hFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000007FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_2}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_11}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFF;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam sdpb_inst_2.INIT_RAM_07 = 256'hFFFFF80000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000003FF;
defparam sdpb_inst_2.INIT_RAM_18 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000;
defparam sdpb_inst_2.INIT_RAM_1A = 256'hFF80000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1C = 256'hFFFFFFFF80000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFC0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000007FFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000007FFFFF;
defparam sdpb_inst_2.INIT_RAM_2B = 256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam sdpb_inst_2.INIT_RAM_2F = 256'hFFFFF80000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_31 = 256'hFFFFFFFFFFF80000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_33 = 256'hF0000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_35 = 256'hFFFFFFE0000000000000000000000000000000000000000FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_37 = 256'hFFFFFFFFFFFFF000000000000000000000000000000000000000007FFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000001FFF;
defparam sdpb_inst_2.INIT_RAM_3A = 256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_3C = 256'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_3E = 256'h00000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_2.INIT_RAM_3F = 256'h037FC7803EF3FFE7BEF9EFFFFFFFDFFFDFFFFC00000000000000000000000000;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_3}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_12}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'h0003FFFFE00000000000001FFFFFFEFFBDFFFFEFDFFF9FFCE7FDFFC5FFF7FBFF;
defparam sdpb_inst_3.INIT_RAM_01 = 256'hF7F9FE007007001CE00FC01E00EFF9CF3F9F3F9FFFFFFFFFFFFFFFFFFFFE0000;
defparam sdpb_inst_3.INIT_RAM_02 = 256'hFF00000003FFFFF000000000000007FFFFFE7F39FE3007DFFF1FF807F8FF807F;
defparam sdpb_inst_3.INIT_RAM_03 = 256'h7F8C3FF3F9FF007007003CF00FC11E00E7F9CF3F8F3F9FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_04 = 256'hFFFFFFFF80000001FFFFFE00000000000001FFFFFE3F1CFE3807CFFF0FF067F8;
defparam sdpb_inst_3.INIT_RAM_05 = 256'hF3E3F87F9F3FF3F9FFE3FFE3F9FCF1FF8F9FFCF3F9CF1F0F3FDFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFFFFFF80000001FFFFFF00000000000001FFFFFF3F9CFE3FE3CFFF0F;
defparam sdpb_inst_3.INIT_RAM_07 = 256'hCFFF07F3F3F87FBF9FF3F8FFF3FFF3F9FCF9FF9F9FFCF3F9E79F0F1FCFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFC0000001FFFFFF800000000000007FFFFF3F9E7E3FE3;
defparam sdpb_inst_3.INIT_RAM_09 = 256'h7E3FF3C7FF27F3F3F83FBF9FFBFCFFF3FFF3F8FE78FF9F8FFE71F9E79F0F9FCF;
defparam sdpb_inst_3.INIT_RAM_0A = 256'h279FCFFFFFFFFFFFFFFFFFFFFFC0000000FFFFFFC00000000000003FFFFF3F9E;
defparam sdpb_inst_3.INIT_RAM_0B = 256'hFF3F9E3E3FF3E7FF27F3F3F9BFFF9FF9FCFFF3FFF3F8FE7CFF9FCFFE79F9E79F;
defparam sdpb_inst_3.INIT_RAM_0C = 256'hF9E79F279FC7FFFFFFFFFFFFFFFFFFFFC0000000FFFFFFE00000000000001FFF;
defparam sdpb_inst_3.INIT_RAM_0D = 256'h000FFFFF1FCF3E3FF3E7FF33F3FBF9BFFF8FF9FCFFF9FFF1FCFE7E7FCFCFFE79;
defparam sdpb_inst_3.INIT_RAM_0E = 256'hCFFE7CF9E3DF279FE7FFFFFFFFFFFFFFFFFFFFC0000000FFFFFFF00000000000;
defparam sdpb_inst_3.INIT_RAM_0F = 256'h0000000007FFFF9FCF3E3FF3E7FF3BFBF9F99FFF8FF9FCFFF9FFF9FCFF3E7FCF;
defparam sdpb_inst_3.INIT_RAM_10 = 256'h3F3FE7CFFE3CF9F3CF27DFE7FFFFE0000000000003FFE00000007FFFFFF80000;
defparam sdpb_inst_3.INIT_RAM_11 = 256'hF800000000000003FFFF9FCF9E3FF1E7FF39F9F9F9CFFF1FF9FCFFF9FFF9FCFF;
defparam sdpb_inst_3.INIT_RAM_12 = 256'h01FCFF3F1FF3C7C03EF9F3CF33CFE7FFFFC0000000000003FFE00000007FFFFF;
defparam sdpb_inst_3.INIT_RAM_13 = 256'h7FFFFFFC00000000000001FFFF9FEF9E3F11E7FF39FC79F9CFFE1FFCFE7FF9FF;
defparam sdpb_inst_3.INIT_RAM_14 = 256'h7FF8FF19FE7F3F8FF007C03E79F3EE73CFE7FFFFE0000000000000FFF0000000;
defparam sdpb_inst_3.INIT_RAM_15 = 256'h0000003FFFFFFE00000000000000FFFF9FE7CE3F11E3FF3DFC10F9C7F83FFCFE;
defparam sdpb_inst_3.INIT_RAM_16 = 256'hFFFCFE7FFCFF18FE7F3FCFF807C33F39F3E673CFE3FFFFE0000000000000FFF0;
defparam sdpb_inst_3.INIT_RAM_17 = 256'h007FF00000003FFFFFFE00000000000000FFFFDFE7CE3F01F3FF3CFE00F9E7F0;
defparam sdpb_inst_3.INIT_RAM_18 = 256'hF8E7E0FFFCFE7FFCFFF8FE7F9FC7F003FF3F39F3E673E7F3FFFFF00000000000;
defparam sdpb_inst_3.INIT_RAM_19 = 256'hE00000007FF80000003FFFFFFF000000000000007FFFCFE7E63FF8F3FF3C7E08;
defparam sdpb_inst_3.INIT_RAM_1A = 256'h007C7CF803E7FFFCFF7FFCFFFCFE7F9FE7F3F3FF1F39F1E673E7F3FFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1B = 256'hFFFFFFF00000003FF80000001FFFFFFF000000000000003FFFCFE7E63FFCF3FF;
defparam sdpb_inst_3.INIT_RAM_1C = 256'hFCF3FF007C7CF803E7FFFC7F3FFCFFFCFF3F9FF3F3F3FF9F99F9E679E7F3FFFF;
defparam sdpb_inst_3.INIT_RAM_1D = 256'hF3FFFFFFFFFFF80000003FF80000001FFFFFFF000000000000001FFFCFE3E63F;
defparam sdpb_inst_3.INIT_RAM_1E = 256'hF3F23FFC79FF1E3C7C78F1E7FFFE7F3FFCFFFCFF3F9FF1F3F3FF9F99F9E279E7;
defparam sdpb_inst_3.INIT_RAM_1F = 256'hF279E3F3FFFFFFFFFFFC0000003FFC0000000FFFFFFF800000000000001FFFE7;
defparam sdpb_inst_3.INIT_RAM_20 = 256'h0FFFE7F3F23FFC79FF3F3E7E78F9E7FBFE7F3FFE7FFC7F3F9FF9F3F3FF9FD9F9;
defparam sdpb_inst_3.INIT_RAM_21 = 256'h9FC1F9F0F9F3F1FFFFFFFFFFFC0000001FFC0000000FFFFFFF80000000000000;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h0000000FFFE7F3F83FFE79F73F9E7E79FCE7FBFE7F3FFE7FFE7F3F8FF8F3F1FF;
defparam sdpb_inst_3.INIT_RAM_23 = 256'hF1F9FF8FE1FCF0FDF3F1FFFFFFFFFFFE0000001FFC0000000FFFFFFF80000000;
defparam sdpb_inst_3.INIT_RAM_24 = 256'h00000000000007FFE3F3F83FFE79E33F9E7E79FCE7F3FF7F1FFE7FFE7F1FCFFC;
defparam sdpb_inst_3.INIT_RAM_25 = 256'h9FCFFE79F9FF8FE1FCF0FCF1F1FFFFFFFFFFFF0000000FFE0000000FFFFFFF80;
defparam sdpb_inst_3.INIT_RAM_26 = 256'hFFFF8000000000000003FFF3F3FC3FFE7CE33FCE7E79FC73F3FF1F1FFE7FFE7F;
defparam sdpb_inst_3.INIT_RAM_27 = 256'h7FFE3F9FCFFE39F9FFCFF1FCF0FCF9F1FFFFFFFFFFFF0000000FFE00000007FF;
defparam sdpb_inst_3.INIT_RAM_28 = 256'h0007FFFFFFC000000000000003FFF1E3FC3FFE3CE33FCE7E39FE71F3FF9F1FFF;
defparam sdpb_inst_3.INIT_RAM_29 = 256'h803FFF7FC03F9FEF8039F9F00FF1FEF9FCFC03FFFFFFFFFFFF8000000FFE0000;
defparam sdpb_inst_3.INIT_RAM_2A = 256'hFF00000003FFFFFFC000000000000001FFF803FE7F803E073FCE7F39FE7803FF;
defparam sdpb_inst_3.INIT_RAM_2B = 256'h7C07FFE07FFF7F803F9FEF0039FDE00FF1FEF9FEFE03FFFFFFFFFFFF80000007;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h000007FF00000003FFFFFFC000000000000001FFFC07FE7F803F07BFE67F39FF;
defparam sdpb_inst_3.INIT_RAM_2D = 256'hFFFFFFFE0FFFE07FFFFFC07FFFFF807FFFF00FFFFEFDFFFF07FFFFFFFFFFFFC0;
defparam sdpb_inst_3.INIT_RAM_2E = 256'hFFFFC0000007FF80000003FFFFFFC000000000000001FFFE0FFFFF807F0FFFFF;
defparam sdpb_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_30 = 256'hFFFFFFFFFFE0000003FF80000001FFFFFFC000000000000000FFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFE0000003FF80000001FFFFFFC000000000000000FFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFE0000003FFC0000001FFFFFFC0000000000000007F;
defparam sdpb_inst_3.INIT_RAM_35 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001FFC0000000FFFFFF800000000000;
defparam sdpb_inst_3.INIT_RAM_37 = 256'h00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001FFC0000000FFFFFF800000;
defparam sdpb_inst_3.INIT_RAM_39 = 256'h80000000000000003FFFFFFFFFFF33FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFC0000000FFFFFF;
defparam sdpb_inst_3.INIT_RAM_3B = 256'h7FFFFF80000000000000003FFFFFFFFFFF23FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFE0000000;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h0000007FFFFF80000000000000001FFFFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFE0;
defparam sdpb_inst_3.INIT_RAM_3F = 256'h00FFF00000007FFFFF00000000000000001FFFFFFFFFFF87FFFFFFFFFFFFFFFF;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_4}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_13}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b0;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000;
defparam sdpb_inst_4.INIT_RAM_01 = 256'hFC0000007FF00000003FFFFF00000000000000001FFFFFFFFFFFC7FFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_03 = 256'hFFFFFFFC0000007FF00000003FFFFF00000000000000001FFFFFFFFFFFC7FFFF;
defparam sdpb_inst_4.INIT_RAM_04 = 256'hCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFE0000007FF80000001FFFFE00000000000000000FFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_06 = 256'hCFCFFF01FFF3F9FFDFEFFE00FF800FFF03FFFC03FF003FF3F7FF007FFFCFFC01;
defparam sdpb_inst_4.INIT_RAM_07 = 256'hCFFC00FFFFFFFFFFFFFE0000003FF80000001FFFFE00000000000000000FF9FF;
defparam sdpb_inst_4.INIT_RAM_08 = 256'h0FF1FF87C7FE00FFE1F0FF8FC7FC007F8007FE00FFF001FE001FE1E1FF003FFF;
defparam sdpb_inst_4.INIT_RAM_09 = 256'h003FFF87FC007FFFFFFFFFFFFE0000003FF80000001FFFFC0000000000000000;
defparam sdpb_inst_4.INIT_RAM_0A = 256'h00000007F0FF8787FE007FE1E0FF87C7FC007F8007FE007FF001FE001FE1E1FF;
defparam sdpb_inst_4.INIT_RAM_0B = 256'hF0E1FF001FFF87FC007FFFFFFFFFFFFE0000001FFC0000000FFFF80000000000;
defparam sdpb_inst_4.INIT_RAM_0C = 256'h00000000000007F0FFC3C7FC003FE1E0FF87C7FE007F8007FC007FF001FF001F;
defparam sdpb_inst_4.INIT_RAM_0D = 256'hFF003FF871FF801FFFC7FC007FFFFFFFFFFFFF0000001FFC0000000FFFF80000;
defparam sdpb_inst_4.INIT_RAM_0E = 256'hF0000000000000000007F8FFE1C7FC183FF1E0FF87C3FF007FC007FC183FF000;
defparam sdpb_inst_4.INIT_RAM_0F = 256'h1FF0F0FFF1FFF831FFFE1FFFC7FFF87FFFFFFFFFFFFF0000001FFC0000000FFF;
defparam sdpb_inst_4.INIT_RAM_10 = 256'h0007FFE0000000000000000003F8FFE0C7FC3C1FF1E0FFC7C3FFFC7FFC7FFC3C;
defparam sdpb_inst_4.INIT_RAM_11 = 256'h7FF87E1FF1F8FFF1FFFC31FFFF1FFFC7FFFC7FFFFFFFFFFFFF8000000FFE0000;
defparam sdpb_inst_4.INIT_RAM_12 = 256'hFE00000007FFC0000000000000000003F8FFF0C7FC7E1FF1C0FFC7C3FFFC3FFC;
defparam sdpb_inst_4.INIT_RAM_13 = 256'hFC3FFC7FF87F1FF1F8FFF1FFFE11FFFF1FFFC7FFFC7FFFFFFFFFFFFF8000000F;
defparam sdpb_inst_4.INIT_RAM_14 = 256'h00000FFE00000007FF80000000000000000003F87FF807FC7F1FF1C07FC7C3FF;
defparam sdpb_inst_4.INIT_RAM_15 = 256'hC0C3FFFC3FFC7FF87F0FF0F8FFF0FFFF01FFFF1FFFC3FFF87FFFFFFFFFFFFF80;
defparam sdpb_inst_4.INIT_RAM_16 = 256'hFFFFC0000007FF00000003FE00000000000000000003F87FFC03FFFF1FF0C07F;
defparam sdpb_inst_4.INIT_RAM_17 = 256'hF0C07FC003FF003FFC7FF87F0FF070FFF0FFFF01FFC01FFFC3FE007FFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_18 = 256'hFFFFFFFFFFC0000007FF00000001F800000000000000000003F87FFC03FFFF0F;
defparam sdpb_inst_4.INIT_RAM_19 = 256'hFFFF0FF0C47FC003FF003FFC3FF87F8FF800FFF8FFFF01FF801FFFC3FE003FFF;
defparam sdpb_inst_4.INIT_RAM_1A = 256'h003FFFFFFFFFFFFFC0000007FF800000000000000000000000000001F87FFC03;
defparam sdpb_inst_4.INIT_RAM_1B = 256'h7FFC03FFFF0FF8847FC003FF003FFC3FF87F8FF800FFF8FFFF00FF801FFFE3FE;
defparam sdpb_inst_4.INIT_RAM_1C = 256'hFFE3FF003FFFFFFFFFFFFFE0000003FF800000000000000000000000000001FC;
defparam sdpb_inst_4.INIT_RAM_1D = 256'h0001FC7FFC03FFFF8FF80C7FC001FF803FFC3FFC7F8FFC00FFF8FFFF00FFC01F;
defparam sdpb_inst_4.INIT_RAM_1E = 256'hFFFF0FFFE3FFFC3FFFFFFFFFFFFFE0000003FF80000000000000000000000000;
defparam sdpb_inst_4.INIT_RAM_1F = 256'h0000000001FC7FF803FFFF8FF80C7FC3E1FFFE1FFE3FFC7F8FFC00FFF8FFFE00;
defparam sdpb_inst_4.INIT_RAM_20 = 256'hFFFE10FFFF0FFFE3FFFE3FFFFFFFFFFFFFE0000003FFC0000000000000000000;
defparam sdpb_inst_4.INIT_RAM_21 = 256'h0000000000000001FC7FF863FFFF8FF80C7FC3E1FFFE1FFE3FFC7F8FF8387FF8;
defparam sdpb_inst_4.INIT_RAM_22 = 256'h787FF8FFFC38FFFF8FFFE3FFFE3FFFFFFFFFFFFFF0000001FFC0000000000000;
defparam sdpb_inst_4.INIT_RAM_23 = 256'h0000000000000000000001FC3FF0E3FE3F8FF81C7FE3F1FFFE1FFE3FFC3F8FF8;
defparam sdpb_inst_4.INIT_RAM_24 = 256'h3F0FF8787FF8FFFC38FFFF8FFFE3FFFE3FFFFFFFFFFFFFF0000001FFC0000000;
defparam sdpb_inst_4.INIT_RAM_25 = 256'h0000007FFFFF0000000000000001FC3FF0E3FE1F0FF81C3FE3F1FFFF1FFE1FFC;
defparam sdpb_inst_4.INIT_RAM_26 = 256'hFE1FFE1F0FF87C7FF87FF838FFFF8FFFE3FFFE3FFFFFFFFFFFFFF8000000FFE0;
defparam sdpb_inst_4.INIT_RAM_27 = 256'h00FFE00000007FFFFF8000000000000001FC3FF0E3FE1F0FF81C3FE3F1FFFE1F;
defparam sdpb_inst_4.INIT_RAM_28 = 256'hFF801FFE1FFE0E0FF87C7FF87FF878FFC00FF801FF003FFFFFFFFFFFFFF80000;
defparam sdpb_inst_4.INIT_RAM_29 = 256'hF8000000FFE00000007FFFFFF000000000000001FE3FE1E1FF060FFC3C3FE3F0;
defparam sdpb_inst_4.INIT_RAM_2A = 256'h3FE3F0FF001FFE1FFF001FF87C7FF87FF8787F8007F001FE003FFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2B = 256'hFFFFFFFC0000007FF00000003FFFFFF800000000000001FE3FE1E1FF001FFC3E;
defparam sdpb_inst_4.INIT_RAM_2C = 256'h1FFC3E3FE3F0FF000FFF1FFF801FF87C3FFC7FF0787F8007F001FE001FFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFFFC0000007FF00000003FFFFFFC00000000000001FE3FE1E1FF80;
defparam sdpb_inst_4.INIT_RAM_2E = 256'hE1FFC03FFC3E3FE1F8FF000FFF1FFFC03FF87C3FFC7FF0F87F8007F001FE001F;
defparam sdpb_inst_4.INIT_RAM_2F = 256'hFF003FFFFFFFFFFFFFFC0000007FF80000001FFFFFFE00000000000001FE3FC3;
defparam sdpb_inst_4.INIT_RAM_30 = 256'hFE3FE3F1FFE03FFC7E3FF3F9FF801FFF1FFFC03FFC7E7FFC7FF0FCFFC00FF801;
defparam sdpb_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC0000003FF80000001FFFFFFF00000000000001;
defparam sdpb_inst_4.INIT_RAM_32 = 256'h000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000003FF80000001FFFFFFF80000000;
defparam sdpb_inst_4.INIT_RAM_34 = 256'h000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000001FFC0000000FFFFFFFC0;
defparam sdpb_inst_4.INIT_RAM_36 = 256'hFFFFC0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001FFC0000000FFF;
defparam sdpb_inst_4.INIT_RAM_38 = 256'h000FFFFFFFE0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001FFC0000;
defparam sdpb_inst_4.INIT_RAM_3A = 256'hFE0000000FFFFFFFE0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000F;
defparam sdpb_inst_4.INIT_RAM_3C = 256'h00000FFE00000007FFFFFFF0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam sdpb_inst_4.INIT_RAM_3E = 256'hFFFF8000000FFE00000007FFFFFFF0000000000001FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_5}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_14}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b0;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'hFFFFFFFFFF80000007FF00000007FFFFFFF8000000000003FFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFC0000007FF00000007FFFFFFF8000000000003FFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFC0000007FF80000007FFFFFFF8000000000003FFFF;
defparam sdpb_inst_5.INIT_RAM_05 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000003FF80000007FFFFFFFC0000000000;
defparam sdpb_inst_5.INIT_RAM_07 = 256'h00000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_08 = 256'h0FFDFDFCF9F9FF9FE01FFFFFFFFFFFFFFFE0000003FF80000007FFFFFFFC0000;
defparam sdpb_inst_5.INIT_RAM_09 = 256'hFC000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07FFFDFDFFFC01F007E0;
defparam sdpb_inst_5.INIT_RAM_0A = 256'hF003C007F8F8F8F0F1FF0FC00FFFFFFFFFFFFFFFE0000003FFC0000003FFFFFF;
defparam sdpb_inst_5.INIT_RAM_0B = 256'hFFFFFFFC000000000003FFE3E3C7E3C00F9FFF87FE007F87FE03FFF8F8FFF800;
defparam sdpb_inst_5.INIT_RAM_0C = 256'h7FF800F003C007F8F8F8F0F1FE0FC00FFFFFFFFFFFFFFFE0000001FFC0000003;
defparam sdpb_inst_5.INIT_RAM_0D = 256'h000003FFFFFFFC000000000007FFE3E3C3E3C00F8FFF87FC007F87FC01FFF8F8;
defparam sdpb_inst_5.INIT_RAM_0E = 256'hFFF8F87FF800F003C007F8F8F8F871FE07E007FFFFFFFFFFFFFFF0000001FFC0;
defparam sdpb_inst_5.INIT_RAM_0F = 256'h00FFE0000003FFFFFFFE000000000007FFE3E1E3E3C00F8FFF83FC007F83FC00;
defparam sdpb_inst_5.INIT_RAM_10 = 256'h83FC30FFF87C7FFC00F001E007F8F8F87C30FE07E007FFFFFFFFFFFFFFF00000;
defparam sdpb_inst_5.INIT_RAM_11 = 256'hF8000000FFE0000003FFFFFFFE000000000007FFE3F1E3E3C00F8FFF83FC007F;
defparam sdpb_inst_5.INIT_RAM_12 = 256'hFC7C7F83FC78FFFC7C7FFF87FFE1FC3FF8F8F87E18FE07FF87FFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_13 = 256'hFFFFFFF8000000FFE0000003FFFFFFFE000000000007FFE1F1E1E3FF8F8FFF81;
defparam sdpb_inst_5.INIT_RAM_14 = 256'h87FF81FC7C7F81FC787FFC7C7FFFC7FFF1FE3FF8F87C7E18FE03FFC7FFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_15 = 256'hFFFFFFFFFFFFF80000007FF0000007FFFFFFFE00000000000FFFF1F1F1E3FF87;
defparam sdpb_inst_5.INIT_RAM_16 = 256'hE3FFC7C7FF81FC7C7F81FEF87FFC7C7FFFC7FFF1FE3FF8787C7F00FE23FFC7FF;
defparam sdpb_inst_5.INIT_RAM_17 = 256'hFFC7FFFFFFFFFFFFFFFC0000007FF0000007FFFFFFFE00000000000FFFF1F1F1;
defparam sdpb_inst_5.INIT_RAM_18 = 256'hF1F1F1E3FFC7C7FF88FC7C3F88FFF87FFC7C3FFFC7FFF1FE3FFC7C7C7F80FE23;
defparam sdpb_inst_5.INIT_RAM_19 = 256'h807E31F807FFFFFFFFFFFFFFFC0000007FF0000007FFFFFFFC00000000000FFF;
defparam sdpb_inst_5.INIT_RAM_1A = 256'h001FFFF1F1F8E3F007C7FF88FC3C3F08FFC07FFC7C3FFFC7FC01FE3FFC7C7C3F;
defparam sdpb_inst_5.INIT_RAM_1B = 256'h7C7C3FC07E31F003FFFFFFFFFFFFFFFC0000003FF8000007FFFFFFFC00000000;
defparam sdpb_inst_5.INIT_RAM_1C = 256'h000000001FFFF1F0F8E3E007C7FF887E003F08FF807FFC3E3FFFC7F801FE3FFC;
defparam sdpb_inst_5.INIT_RAM_1D = 256'hFE1FFC3C3E3F807E31F003FFFFFFFFFFFFFFFE0000003FF8000007FFFFFFFC00;
defparam sdpb_inst_5.INIT_RAM_1E = 256'hFFFC00000000001FFFF1F8F863E007C7FF0C7E003F1C7F00FFFC3E3FFFC3FC01;
defparam sdpb_inst_5.INIT_RAM_1F = 256'hC3FC00FF1FFC3E3E3F807E38F803FFFFFFFFFFFFFFFE0000003FF8000007FFFF;
defparam sdpb_inst_5.INIT_RAM_20 = 256'h0FFFFFFFF800000000003FFFF0F8FC67F007C7FF0C7F003F1C7E01FFFE3E3FFF;
defparam sdpb_inst_5.INIT_RAM_21 = 256'h3E3FFFE3FEE0FF1FFE3E3E3F807E38F803FFFFFFFFFFFFFFFE0000001FF00000;
defparam sdpb_inst_5.INIT_RAM_22 = 256'hF000000FFFFFFFF800000000003FFFF8F8FC47F803C3FF0C3F003F0C7E03FFFE;
defparam sdpb_inst_5.INIT_RAM_23 = 256'h1FFFFE3E1FFFE3FFF8FF1FFE3E3E3F0C7E007FE3FFFFFFFFFFFFFFFF0000001F;
defparam sdpb_inst_5.INIT_RAM_24 = 256'h00000FF000000FFFFFFFF800000000007FFFF8F8FE07FFC3E39F003F0E1F003E;
defparam sdpb_inst_5.INIT_RAM_25 = 256'h1F003E1FFFFE1F1FFFE3FFF8FF1FFE3E3E3F0C3E007FE3FFFFFFFFFFFFFFFF00;
defparam sdpb_inst_5.INIT_RAM_26 = 256'h0000000000000000001FFFFFFFF000000000007FFFF8F87E07FFE3E38F003F0E;
defparam sdpb_inst_5.INIT_RAM_27 = 256'h001F1F1F001E3F3FFF1F1FFFE1FFF8FF1FFE3E3E3F1E3E007FE3FFFFFFFFFF80;
defparam sdpb_inst_5.INIT_RAM_28 = 256'hFFFF800000000000000000001FFFFFFFF00000000000FFFFF8787E07FFE3E38F;
defparam sdpb_inst_5.INIT_RAM_29 = 256'hE3E38F001F1F1F001E3E1FFF1F1FFFE1FFF8FF1FFE3E1E3F1E3E003FE1FFFFFF;
defparam sdpb_inst_5.INIT_RAM_2A = 256'hFFFFFFFFFF800000000000000000003FFFFFFFE00000000001FFFFF8787F07FF;
defparam sdpb_inst_5.INIT_RAM_2B = 256'h7F07FBE3E18F000F1F1F000E1C1FFF0E1FFFF1FE00FF0FC01F0C3E1E3E003FE1;
defparam sdpb_inst_5.INIT_RAM_2C = 256'h3E3FF1FFFFFFFFFF800000000000000000007FFFFFFFC00000000001FFFFFC38;
defparam sdpb_inst_5.INIT_RAM_2D = 256'hFFFC107F07F003E10F1F8F0F0F1F0F0C1FFF801FFFF1FC007F0F801F003E1E3C;
defparam sdpb_inst_5.INIT_RAM_2E = 256'h3E1E3C3E1FF1FFFFFFFFFF80000000000000000000FFFFFFFF800000000003FF;
defparam sdpb_inst_5.INIT_RAM_2F = 256'h0007FFFFFE00FF87F001F00F1F8F0F0E1F8F003FFF801FFFF1FC007F8F801F00;
defparam sdpb_inst_5.INIT_RAM_30 = 256'h801F803C3E3C3F1FF1FFFFFFFFFFFFFFFFC0000007FFFFFFFFFFFFFF00000000;
defparam sdpb_inst_5.INIT_RAM_31 = 256'h000000000FFFFFFE00FF87F001F00E1F870F8E1F87803FFFC03FFFF1FC007F8F;
defparam sdpb_inst_5.INIT_RAM_32 = 256'h007F8F801FC07E3F3E7F1FF9FFFFFFFFFFFFFFFFE0000003FFFFFFFFFFFFFE00;
defparam sdpb_inst_5.INIT_RAM_33 = 256'hFFF800000000001FFFFFFF01FFC7F001F81F1FC79F9F3F8F807FFFC07FFFF1FE;
defparam sdpb_inst_5.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000003FFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_35 = 256'hFFFFFFFFE000000000003FFFFFFFC3FFFFFFFFFE3FFFFFFFFFFFFFF1FFFFF8FF;
defparam sdpb_inst_5.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000001FFFF;
defparam sdpb_inst_5.INIT_RAM_37 = 256'h00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000;
defparam sdpb_inst_5.INIT_RAM_39 = 256'hF0000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3B = 256'hFFFFFFF0000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3D = 256'hFFFFFFFFFFFFF800000000000000000000000000001FFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFF800000000000000000000000000003FFFFFFFFFFFFFFF;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_6}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_15}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b0;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000003FFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000001FFFFF;
defparam sdpb_inst_6.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000003FFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000003FFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000001F;
defparam sdpb_inst_6.INIT_RAM_0C = 256'h00001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam sdpb_inst_6.INIT_RAM_0E = 256'hFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_10 = 256'hFFFFFFFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000003FFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000003FFFF;
defparam sdpb_inst_6.INIT_RAM_1F = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000;
defparam sdpb_inst_6.INIT_RAM_21 = 256'hE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_23 = 256'hFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_25 = 256'hFFFFFFFFFFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFF;
defparam sdpb_inst_6.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000003F;
defparam sdpb_inst_6.INIT_RAM_34 = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00;
defparam sdpb_inst_6.INIT_RAM_36 = 256'hFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_38 = 256'hFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_6.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_7}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_16}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b0;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFF;
defparam sdpb_inst_7.INIT_RAM_07 = 256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam sdpb_inst_7.INIT_RAM_09 = 256'hE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0B = 256'hFFFFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0D = 256'hFFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000007FFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007F;
defparam sdpb_inst_7.INIT_RAM_1C = 256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_7.INIT_RAM_1E = 256'hFFFE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_20 = 256'hFFFFFFFFFE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007FFFF;
defparam sdpb_inst_7.INIT_RAM_2F = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000;
defparam sdpb_inst_7.INIT_RAM_31 = 256'hC0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_33 = 256'hFFFFFFE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_35 = 256'hFFFFFFFFFFFFE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFE0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000FFFFFFFFFFFFFF;

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[30:0],sdpb_inst_8_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_8}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_17}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_8.READ_MODE = 1'b0;
defparam sdpb_inst_8.BIT_WIDTH_0 = 1;
defparam sdpb_inst_8.BIT_WIDTH_1 = 1;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_8.RESET_MODE = "SYNC";
defparam sdpb_inst_8.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000007F;
defparam sdpb_inst_8.INIT_RAM_04 = 256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sdpb_inst_8.INIT_RAM_06 = 256'hFFFE0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_08 = 256'hFFFFFFFFFE0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFF0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000001FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000FFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000FFFFF;
defparam sdpb_inst_8.INIT_RAM_17 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000;
defparam sdpb_inst_8.INIT_RAM_19 = 256'hF0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1B = 256'hFFFFFFF8000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1D = 256'hFFFFFFFFFFFFF8000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFC000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000001FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000001FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000FFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000FFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000FF;
defparam sdpb_inst_8.INIT_RAM_2C = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam sdpb_inst_8.INIT_RAM_2E = 256'hFFFFF800007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_30 = 256'hFFFFFFFFFFFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0001FFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003FFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_8.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF803FFFFF;
defparam sdpb_inst_8.INIT_RAM_3F = 256'h00000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[17]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[16]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[15]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(sdpb_inst_2_dout[0]),
  .I1(sdpb_inst_3_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(sdpb_inst_4_dout[0]),
  .I1(sdpb_inst_5_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(sdpb_inst_6_dout[0]),
  .I1(sdpb_inst_7_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_2)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_2)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_5),
  .I1(mux_o_6),
  .S0(dff_q_1)
);
MUX2 mux_inst_10 (
  .O(dout[0]),
  .I0(mux_o_8),
  .I1(sdpb_inst_8_dout[0]),
  .S0(dff_q_0)
);
endmodule //Gowin_SDPB4
