//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.10
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Wed Sep 06 14:26:27 2023

module Gowin_SDPB5 (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);//sobel_3x3_v2

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [14:0] ada;
input [7:0] din;
input [14:0] adb;

wire lut_f_0;
wire lut_f_1;
wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [1:1] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [2:2] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [3:3] sdpb_inst_3_dout;
wire [30:0] sdpb_inst_4_dout_w;
wire [4:4] sdpb_inst_4_dout;
wire [30:0] sdpb_inst_5_dout_w;
wire [5:5] sdpb_inst_5_dout;
wire [30:0] sdpb_inst_6_dout_w;
wire [6:6] sdpb_inst_6_dout;
wire [30:0] sdpb_inst_7_dout_w;
wire [7:7] sdpb_inst_7_dout;
wire [29:0] sdpb_inst_8_dout_w;
wire [1:0] sdpb_inst_8_dout;
wire [29:0] sdpb_inst_9_dout_w;
wire [3:2] sdpb_inst_9_dout;
wire [29:0] sdpb_inst_10_dout_w;
wire [5:4] sdpb_inst_10_dout;
wire [29:0] sdpb_inst_11_dout_w;
wire [7:6] sdpb_inst_11_dout;
wire [27:0] sdpb_inst_12_dout_w;
wire [3:0] sdpb_inst_12_dout;
wire [27:0] sdpb_inst_13_dout_w;
wire [7:4] sdpb_inst_13_dout;
wire [23:0] sdpb_inst_14_dout_w;
wire [7:0] sdpb_inst_14_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire mux_o_6;
wire mux_o_8;
wire mux_o_16;
wire mux_o_18;
wire mux_o_26;
wire mux_o_28;
wire mux_o_36;
wire mux_o_38;
wire mux_o_46;
wire mux_o_48;
wire mux_o_56;
wire mux_o_58;
wire mux_o_66;
wire mux_o_68;
wire mux_o_76;
wire mux_o_78;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ada[11]),
  .I1(ada[12]),
  .I2(ada[13]),
  .I3(ada[14])
);
defparam lut_inst_0.INIT = 16'h4000;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(adb[11]),
  .I1(adb[12]),
  .I2(adb[13]),
  .I3(adb[14])
);
defparam lut_inst_1.INIT = 16'h4000;
SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b1;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h263D3F59F81D5E8E63684C3ED6BFCCD90EC5417E27FAF4FE5AEE4F1BA7D60F34;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h10777B6F5E067763FA766D0049BF7432079290021C7F729E5CDBF5FF5B3DE7A6;
defparam sdpb_inst_0.INIT_RAM_02 = 256'hC904102CABDC36492A31B7F7A0E54E415D3A2EEE17DC3C30706CEE4AD7462058;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h01093BE42C40A842082523EC1FEAC146CEDF3B9F908CDE3F5FEF4330848CAF85;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h05111F2BD4F3003082110FA0CB6300F6D149EF263FB1BC935AF43F8E0B7D200E;
defparam sdpb_inst_0.INIT_RAM_05 = 256'hB3A7633F21E20E1273DA45AE28380FE7A97851F91F65587D5D4E1CB94964FF5B;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h8C6C13DFF831F599FF39A760BA8270D5F44E03355322A18FDC9046E2F5B20696;
defparam sdpb_inst_0.INIT_RAM_07 = 256'hF326783FBE302FFB89A099B82F086CCFF6F3D6B7D2C30CB3BE90401639F936BD;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h0AC09CDEFD5C128DAD5BA2DB4880EF7C3F15944F9BA3057D3F60C9D0C85BB62D;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h1C7E2200C0880E15397F00DCF178428D1840B8478348167F41641BA70B9C0889;
defparam sdpb_inst_0.INIT_RAM_0A = 256'hEEDF194501730F076F4410140787BFAB4CFFBD03BA843F91DAA819796F477C01;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h78876C55DE6DE9765F2E83E3D168A40193BCFF91F7834B518E50B7D5EAF7D04C;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h5F2CE7856C61D2CF0D04445B0F52D38278EC6F8048FAEBE2849572868B355BF0;
defparam sdpb_inst_0.INIT_RAM_0D = 256'hAA74D6D53B475258D54EFF48FE4A53E791DE053283D937A7107F1CF6E64AC7DE;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h8E11E39D6A77EF07879F6EEF7BF252A16B3258872C9BC94FEA2F0CCFA86AF6DE;
defparam sdpb_inst_0.INIT_RAM_0F = 256'hDDF89AD386B00BF074CFDB0675A9902D1773A3DEF22B691BF5E6330FD3272268;
defparam sdpb_inst_0.INIT_RAM_10 = 256'hA5CE65F801C40726C961802B9F47FB45A0A133B69699F0134A41C0744D8ED14A;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h12B765CA9B2B4F5363A077FB90427812FABE762FF3853D1F3096D4C4908AFB22;
defparam sdpb_inst_0.INIT_RAM_12 = 256'hE02D0DBB7DE96B86A3BCC19B602F307F3C3A961D5FAED1B6E5F0900EB1A5D912;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h42F88137FE503FF7F8541C2C36F14267FBF6D807817BFD542FAC56C111D8BC65;
defparam sdpb_inst_0.INIT_RAM_14 = 256'hF0F6F19FBD0D8D05BD4A03FFB17D56C349916C96CDE134E4356F452BCA6BBA67;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h2ACF9FEF82FF7DA3356F3B17C9A40329DEAFFC2E5F79056D13AA46F64EADABF6;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h2490ED363D7369E9B44BCBBEA7B61CED3F7FAA3FF2E24FD8A193467530AB158D;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h07F4CCF750CA2172FE9E6D66DE077E9F99FEAEBC0FE7A3A06A37C7492CB7C784;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h8D841AA1858A71EB5A3A3B7BC340B116BD01ADF9E42A0CF80D5E1E3F369A70BD;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h513FE72FAB5DC7752167897E74E1E4956D8693D35B06FFFDE43F7C3B959AE556;
defparam sdpb_inst_0.INIT_RAM_1A = 256'hDFF3B1A3EA9A9CDA4D47875F070A25BDA02213933974766BF52877F5BA1D24E2;
defparam sdpb_inst_0.INIT_RAM_1B = 256'hA4D552FE7FD112D746FFA21C848CE41DBBCC91B30411785FDE8D5CFA034007FB;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h6C023B32CB211FD6BE218B5E7261891D5BCC9F8D514B9B40C9E04A380A43B60D;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h22B67AFF23C65654B7510ADFB8525579DBA85F921666F89D95AF2C6FE4548C45;
defparam sdpb_inst_0.INIT_RAM_1E = 256'hE0536E169736B354DF1511A771139C3EFD06544C740CB003C5A7E32B8DE1357C;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h9A566E27F2DE4A3BFEA8696227C09C25C5EFF06235FFDFC9245E90D1C4F2B447;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h8893987B23FCCB2FF25C807D01C088DB774874584A85F8719E7F86E9378F47E5;
defparam sdpb_inst_0.INIT_RAM_21 = 256'hF69776E5ABC71FE949D5FB4E99A9B01C5F0098E23025E79F9CF5D020E5AF827C;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h6EE4E78C3EBB4494B517076CBCF0905CD6CAA21893EC4F41A5AFF0B8F890F0B2;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h26B18E26462E2680379E2DCA426BD0A2DBE883B4E540F42AFA9B01DE75438959;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h0CAA8FDB7061A3748F92B8DC2028D489A57E6DA72EFE680A244BE8442614BD62;
defparam sdpb_inst_0.INIT_RAM_25 = 256'hF77D2DBF7A302211ECD9C5F576E228D1888681DEB6FCF15D1D36D90E28E73D59;
defparam sdpb_inst_0.INIT_RAM_26 = 256'hF35708EB7071C3F46FEFF564BA9F492C457D5D00490511F9D7B11C053D61B875;
defparam sdpb_inst_0.INIT_RAM_27 = 256'hDCC07754EAE91E575829584FEB530141017909648E0E39F5583F02F5F7BBE5AB;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h94A27245D8D025CE1910301AF4D6FEF47AFFDAF8D0954850B74F35CA0CE5F377;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h1A37F4310714F033FC3F0158DB8F1A6DED0CD9FA576DE3D5D40483F020A7E976;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h6B0453DA0A39B1829C732B0FFBD2B081249DDC0391E8803DF8D1C8FF55326293;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h16EB44381A0B03F2F74DFFECB296A8261EF3C10EADFFAC30119581A94B6FB32F;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h821280728AAFF912D30E54EDDC1B8F7C857DB08D3EF7775CBA062F6CB2924DD0;
defparam sdpb_inst_0.INIT_RAM_2D = 256'hFFA0913735D710DEA7F67F201C0A80DBFB82F63FB7C828AC5086F970C2D6DE01;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h8D9DEF1F56B27F85005D414848A8BC7C5616E801B8B6724F62B4E0E2807FE318;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h9EA6DADD4483DBE69A798E9E26251CA3A7466128B10F548339FFA277F43838F8;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h4265D45E8F9C5C1F4018BEBDADCC0790EDC37D7B1100A000FA47F1010EBDB060;
defparam sdpb_inst_0.INIT_RAM_31 = 256'hAC1B7BB1F4BA96FEFC0501AB3C50BBFE972592C046F3816EC8B6389C9581ECC6;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h07FBC35C0B032E08BF0A8AC01DD00AC7334D6A77CB5C86A063C7A8F4B1F14DB1;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h27DF31E379119BE23306280172EE38341D0A7071FA23205D5EF5B23C3F2B5D7C;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h714AFB3F0448EE3BE6F99272D126F5022BA40B0B919F8A7A45469B464C77BCA1;
defparam sdpb_inst_0.INIT_RAM_35 = 256'hB74B8E51683FE67CF6465ED37E613C4403E4FB2673517A6506318053F7155BF2;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h8B7852FDDE58CE1F383EC5F6607A20C8878EB0812C487F7E32868A5C9A6049EC;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h04721D10E0CCD1F7DDD6E5C191F7E39D7A189B39EDD2BE4C8E349BF6A44C127D;
defparam sdpb_inst_0.INIT_RAM_38 = 256'hF859AAEA9ABEF2373B70E5F6E3D14673777AEFD1065BC0B21F18620E9D9060F4;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h6001097BBC2261299E9FBF4A480485FD22CA79CC6CE465F4AE46FF5A905EA0C1;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h4FAE01784024A4520DCF276E691B9DF4BE4404FF7593D080F64DAFD3681E3945;
defparam sdpb_inst_0.INIT_RAM_3B = 256'hDC0EFE6DFAD102D8181748BB1E61ABF1FF9E7D208DC4DD7FF7C80F831E5613E7;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h3B9E5B47590D67E030F1D3B2000943A569FA3BA04FD60D2F487767CFFC3C57A5;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h4C9DCF4CBFEFC3406E36ACA06925808E18DBF6C78D46003A6C7B80C5C4BF9863;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h99293648B65CE12AC011B69FFE30E928961C93296CB00978C027C03C62FC3EE4;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h772860080905B02807ACDB9CF042C5E9754B9F14FCA2D172BB8FF830977DF84B;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b1;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h02FFD69E7F9902159EF033FF800027200FFFFFFFFFDEDCFE5FFF901BBFCFF1BA;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h10777F90A006F7F3C77C4C00127F03FE00032FFC1C7FFFFB7EFBF77F5BFF1800;
defparam sdpb_inst_1.INIT_RAM_02 = 256'hE90000042BDC3776D54115FCBBE41000AFDA01FE0004B3CF806CEEDBFF460058;
defparam sdpb_inst_1.INIT_RAM_03 = 256'hFE813BE42C000A00082523F3E0105047E7FC85206FEC21FF400375CF700DAF85;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h0001AF852A0101B082104003000301FD6EB680C67090404CAFFC007F00017F11;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h4877629D80853D07F00245BE28300000407871F9FAB8A00D1BDC4004A7F6013F;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h043C048007DBF027FE033BFE770070DFF440021AA00A21A7FF7FA80235AA0108;
defparam sdpb_inst_1.INIT_RAM_07 = 256'hF7FFFFC840018001D45C9027FE001FF37E83F6B7FEC30080024080165FFFDD42;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h0840201EFFFFFFFC0030000277FFFB43DF10FF4106AD7FFFFF6000505000100D;
defparam sdpb_inst_1.INIT_RAM_09 = 256'hF7FE0000C0800005397FFFFF3C838200A7BFF8003DC84AEC0A786CFFF7FC2008;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h3862933AFFFB0007E54018100FDFEFDFFBC04090453FBF8027E83DF088F47E7E;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h447F2FF5C1B8C94821DE8202D520000013FDFFFF7EFCA46E532FFFC001FFFFFD;
defparam sdpb_inst_1.INIT_RAM_0C = 256'hA0F57F84409FCA7F11FCDE2600BDC032552C000000FEFFFFEFCE894154FABFF0;
defparam sdpb_inst_1.INIT_RAM_0D = 256'hBFFFEF4AC0AEFC580065FE4DC76ECC71B001F44C34F0A000007F1DF6FFFD7821;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h4001E39DFE72FEF84861B7EF0109FD99F4CD206429D831107F9ECC20004AFFFE;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h0FE36CF668880DF6F6DFFFF98A167FFD14C01DA4E650D602D23C0F0010CF6507;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h5BBE1C7801B03D621664082BBF5FFBBADE1ECD7281040FEF531515042E81D3C0;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h52B122C92F08C33340B270D2C5801012FEBF7FFFDC7CC6FF308023FAE4446A58;
defparam sdpb_inst_1.INIT_RAM_12 = 256'hA01402449BE4FBDC6123D8876029FE20D540809D5FFCF1FFFE072FFFB18002ED;
defparam sdpb_inst_1.INIT_RAM_13 = 256'hC6D53EFFFE4000080443859A1C715920FBFF56C3C70400103FBCD6C1B1E503FD;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h50F6F1D7BD1E63FFFF48100041DAA1F4EC074D4E3FFEC19F43209A01CA6BBA77;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h1B27801002FFFFA337FFA4EDF9A4021004DBDDE5E11684330823E04F1BD45409;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h1ED24606BDD25834004BEFFEBFBFA792FF7FAA0000F1335AC4D82EE4F0C07688;
defparam sdpb_inst_1.INIT_RAM_17 = 256'hD038F75FCF16BB6022CB635900077EDFD9FFF153FFE7A3A0003BFF901A4360CA;
defparam sdpb_inst_1.INIT_RAM_18 = 256'hB48723213B7696A6B9DA99C9308032704201FFF9A43BF607F7DE3EFF029C7D95;
defparam sdpb_inst_1.INIT_RAM_19 = 256'hBAFFFFF9685FDFA7B71FECEE2C0AE363AEE6ABF70006FFFFE43FFD84EBFEE7FE;
defparam sdpb_inst_1.INIT_RAM_1A = 256'hFFF3B5BC1FFFFAF16935F5A7E7CA3F18B70080FC135BBF2D350877FF1A153591;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h4F3553FFFFD113D8191FF5DB110799989C172C433D80C34F8F1A6602D14007FF;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h12533F6152691FD7FE61AB57A19FFFE3B6F480C7B57A1F27DA90D1B40D454EBA;
defparam sdpb_inst_1.INIT_RAM_1D = 256'hA099F6C68C0CBAC717DFB7FFF956557B98F7F3EA5C5E4F2EE4B1C78509FCE2BB;
defparam sdpb_inst_1.INIT_RAM_1E = 256'hCB525AB702477C7DB0E82315E6C85EFFDDC6545E2C33FFFC80BC98917B72DF58;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h648782354FCE99B38762DFA10C3FE3AB5B78015DFFFFDFC9BA01EF2E06BEF34A;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h8F7007845C188824A93C311BFBD6A6F68337A0DB609204007EFF86C9BD05B85B;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h31F7F6E7BAA700169003E0287557B3BADE4ACBF8394A0E76CCF8242E4BFFE07C;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h7D4540040A1FC494B119809B0280A1FF9C9297A290AB46C0EDB007AE36040001;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h2C60F0308F4210002E41EFCE427C708C00400285BEAE6916BA51AB3E65C38F63;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h7A7E7D4749C49D3728B95822065B7DBFE579BC1080126FD5E2701C6E9E8D6ADE;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h1BAF4781B0DB6D37C1495C5BDC08DD404F4A7FFCB4FEC711E026DF9519B28BF6;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h1C135F0EAD6B429F89FCACDBB16A6FAF6C36C1140EB68FF9F5B9918084003F9A;
defparam sdpb_inst_1.INIT_RAM_27 = 256'hDDC03F8C01081784D04AE85C0A4910CCC0054FADFF3C637E7FF521F5F7BBBEFC;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h78A6813FF8D027E204A031E31D31F60DBE75BEC4702E9095963FDB08DD6748F7;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h570FFE779E4432AFFC3101FDC010135193C52EBED11C1C2E3C1BFA2D7D9FF331;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h9E0BFBDC1187B3CF9E4559A0FFF2B0C66020003C241BF4B1E7F030FF2D0DFF54;
defparam sdpb_inst_1.INIT_RAM_2B = 256'hD1E4BFC7FA04FFF2F8027FF19FE398BFFEF3C38F1B40043F5DFCFBF1E7E04CC0;
defparam sdpb_inst_1.INIT_RAM_2C = 256'hBC381AE3E9C1FFFFF700AFEDD0007F7F2F51A8B536F677F8C700C029C3765CFB;
defparam sdpb_inst_1.INIT_RAM_2D = 256'hFE1322033E1845AC3601FBFFFC057F7FE90025BFE34CC1238FA1F5E0FDC02001;
defparam sdpb_inst_1.INIT_RAM_2E = 256'hD3FDFF9E565E41053FE194C9EA267F7DD60007FFB8B63EEFF8D80B11C9FFEFB8;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h7FF85DD40BBFFFE6DFE7C90B3FDA1B5BFC229128F1002B7FF9FEAA83FFDB2993;
defparam sdpb_inst_1.INIT_RAM_30 = 256'hFD9125AA7FF3A0419CB3EFFDADF9C200EDFD8193A8B0C880FA000EFFFEFE021F;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h3E86000208E5027E03FEFE0FD94AFBF6F2BE7D0046FFFE2CF0FA33A0DC800109;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h8641775E0E02A000B05E23C0022FFFF81F90A77FFB5F5F2043DFBEC8C1441170;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h26EEF1F7E58CA90E000610016C61CFFC02620FFE132128DFFFF5C7941F2F559F;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h77DEFC0E055AE63BF168EDB9D1E7F1026B63F7F4FDB999FFB827567FFDF7B1E1;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hFFB7501D9E7FE78761445EE37F8BB446E3E0FA67E6C0006158A4153FF8ACA715;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h64A1C35FFFF7E0C527FEC6C1E07E20C987F413BF5C487F3F48448CFF4D16E3DF;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h3BF26C028FB7F46DFFFFEFCA1C7DE7F0BA1C933AEFFF68F31EA41FEE6CCC1E0D;
defparam sdpb_inst_1.INIT_RAM_38 = 256'hDBF9A2E4F0FED35E04E0AF0147DBF8724C87FFFE7E4A603201164C96E790A0D7;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h4003C7ADEDF26426E25FD65A0FFE0FD1C57BFE0BD36BA67B12407F5A005F2E8B;
defparam sdpb_inst_1.INIT_RAM_3A = 256'hF2622161C025D44F947F27DC6A7BE88C01B9D8008997FF7484705FDE0BA81D40;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h1E3A69FDFC3900980807E3781017BBEA0BBEDC88801A5D0008ECEFFCB72FCF6F;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h04604AB8A2D6241F734F93B20009FF6320C7FBFF83CFF61F400036C003CB8FFA;
defparam sdpb_inst_1.INIT_RAM_3D = 256'hCC002EDC80101AFF905E8BEDFE43818E9EDBF8BB22CDFFBF9EA7F5BF84000C60;
defparam sdpb_inst_1.INIT_RAM_3E = 256'hE3C8C9B7FE40033FC00E47A0003BA9EC6FE45A297CA03E580EA07EFFA15BC69F;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h24D49FFFF45C02D7FFEC4319F0001148880A267927DCBB02D7FFFBAA97EC077F;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b1;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'hFD00001F1F990204000FFFFE800000000FFFFFFFFFFEDCFE5FFFFFE4402001B8;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h10777FFFFFF90803FFFC4C000000FFFE000080001C7FFFFFFEFBF7FF5BFFFFFF;
defparam sdpb_inst_2.INIT_RAM_02 = 256'hE90000042BDC377FFFFEEA00BBE400000005FFFE00075000006CEEDBFF460058;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h00013BE42C000800082523FFFFFFAFB847FC01000013FFFF40038800000DAF85;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h0001D079000101B082100000000301FFFFFF7FF980F000000003FFFF000180C0;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h00089FFF808165E2000245BE28300000007871F9FFFFFFF2E45C00000009FFFF;
defparam sdpb_inst_2.INIT_RAM_06 = 256'hFBC0008000040FFFFE034111010070DFF4400210000221AFFFFFFFFDCA420000;
defparam sdpb_inst_2.INIT_RAM_07 = 256'hF7FFFFFFFFFE000000036FDFFE00E03D814FF6B7FEC30080020000167FFFFFFF;
defparam sdpb_inst_2.INIT_RAM_08 = 256'h0840001EFFFFFFFFFFEFC002400004BFFF1080B8D8727FFFFF6000505000100D;
defparam sdpb_inst_2.INIT_RAM_09 = 256'hFFFE0000C0800005397FFFFFFFFFFA00000007FFFFC87518259387FFFFFC0008;
defparam sdpb_inst_2.INIT_RAM_0A = 256'h77ADECBFFFFB0007E74018100FDFFFFFFFFFFEA00000407FFFE8070C731181FF;
defparam sdpb_inst_2.INIT_RAM_0B = 256'hBFFF700C7FD26E85FFFE8203AA20000013FDFFFFFFFFFFC00280003FFFFFF005;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h0000007BBFFFD901C9F8FDE77FFFC003126C000000FEFFFFEFDFFFE00000000F;
defparam sdpb_inst_2.INIT_RAM_0D = 256'hBFFFFFBE000001A7FFFFFBB2857A3F156FFFF400840C2000007F1DF6FFFFFFF8;
defparam sdpb_inst_2.INIT_RAM_0E = 256'h0001E39DFE73FFFF80000010FEFFFF6EBFA07FFAD227F90043083C00004AFFFE;
defparam sdpb_inst_2.INIT_RAM_0F = 256'h0E23F33200800DF6F6DFFFFFE0000002EBBFFFFFDDF02FFC8E03FF001E0F6500;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h18BE03F801C7FB5E0064002BBF5FFBFFF800008D7FFFFFF0BCFC897EA1002FC0;
defparam sdpb_inst_2.INIT_RAM_11 = 256'hEC5F8FE088F7C0F340BA5843C0001012FEBF7FFFFE040000CF7FFFFF02FE6AFE;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h5FFBFFFFEC0E3FFAA01E387F602EABA8F400801D5FFEF1FFFF8000004E7FFFFF;
defparam sdpb_inst_2.INIT_RAM_13 = 256'hC6F8000001BFFFFFFA9015FE542AC71FFBFF8D00330000103FBCD6C1B1E00002;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h50F6F1D7BD1E000000B7FFFFFE0201F7383CBCC1FFFFFB5331E00001CA6BBA77;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h2A93800002FFFFA337FF8000065BFDFFFB37400FE3887B10FFC1DF4B9E8C0000;
defparam sdpb_inst_2.INIT_RAM_16 = 256'h0109B358C24D3800004BEFFEBFBFE080008055FFFF062037DC871E2C0F05257E;
defparam sdpb_inst_2.INIT_RAM_17 = 256'hC013136AC017FC493E55474000077EDFD9FFF80000185C5FFFC308588639BEDA;
defparam sdpb_inst_2.INIT_RAM_18 = 256'h5B783A9CBF010C6B7815276BA3F3DEF00001FFF9A43BFE000021C100FD60237D;
defparam sdpb_inst_2.INIT_RAM_19 = 256'h0400001A0D201984270017B99C0CC0F290E4BCEF0006FFFFE43FFD8000011801;
defparam sdpb_inst_2.INIT_RAM_1A = 256'hFFF3B5B80000000754CE86DC19C8B8FC8F02F37E06DD4CECF50877FF3A1535E0;
defparam sdpb_inst_2.INIT_RAM_1B = 256'h103553FFFFD113DE00000801FE1171C8C2A69AE733817880125F2FF44F4007FF;
defparam sdpb_inst_2.INIT_RAM_1C = 256'hFF882E5C479A9FD7FE61AB5FA000000D000340F5EEC101CDE270BA13F111E5F0;
defparam sdpb_inst_2.INIT_RAM_1D = 256'hCA37FACA7FF55AE02D7F6FFFF956557BF800000247E49A307871286BA54CE278;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h98B5084FFD2CFE6A8FFEF3916E2878FFFDC6545E7C00000070D93C1D8FE81089;
defparam sdpb_inst_2.INIT_RAM_1F = 256'h00200FF66AD6300BBC163F9623FF34437D78037FFFFFDFC9BE00000012D3320C;
defparam sdpb_inst_2.INIT_RAM_20 = 256'h8FF0000000070FDF3259113D4B4D9EED48FFCD7011D00067FEFF86C9BF840000;
defparam sdpb_inst_2.INIT_RAM_21 = 256'h4FF7F6E7BAFF00000000837799986E2FA2A647FCAD3FF7C81958002D3FFFE07C;
defparam sdpb_inst_2.INIT_RAM_22 = 256'hA196C00409FFC494B11F80000080B883B8E37F0A2DDB21C1716FFAF8877C0001;
defparam sdpb_inst_2.INIT_RAM_23 = 256'h29958179C05610003B3FEFCE427FF080004002FA64F06112A51898FE4258716D;
defparam sdpb_inst_2.INIT_RAM_24 = 256'h8CD6E33F411C3F596B5300000707FDBFE579DC0000126F6B35000399810CE63E;
defparam sdpb_inst_2.INIT_RAM_25 = 256'h25032381DB1EE30FC06A6F0ACDF394400F69FFFCB4FEFF100026DFF1921D87FF;
defparam sdpb_inst_2.INIT_RAM_26 = 256'h00135FF26B8D29800DB863C7B00E5516F8F8F8840F8E7FF9F5B99F8004003FE1;
defparam sdpb_inst_2.INIT_RAM_27 = 256'hDDC03FFC000817F89F57D2C3F4580FC3C001D1D1F2FFA19CFFC59FF5F7BBBF7C;
defparam sdpb_inst_2.INIT_RAM_28 = 256'h1D4968FFF8D027FE000031FC3B0F78A3FEF32EC3F00011FB72FFE7F2001467F7;
defparam sdpb_inst_2.INIT_RAM_29 = 256'h6EFFFFAFE9D44E5FFC3101FFC000137E18AA4129D103E001FC000358647FFDEE;
defparam sdpb_inst_2.INIT_RAM_2A = 256'hFE0004201F7FB3F5BC0CC71FFFF2B0C7E000003FC69B80A4600FFF00FD000018;
defparam sdpb_inst_2.INIT_RAM_2B = 256'hB01FFFFFFA00000D007FFFFECD208651FEF3C38FFB40043FE12EC583201FFFFF;
defparam sdpb_inst_2.INIT_RAM_2C = 256'hBFDCB7CF583FFFFFF70000122FFFFF7FCA314774FEF677F8FF000029FC671662;
defparam sdpb_inst_2.INIT_RAM_2D = 256'hFFF200033FE09CA56E0FFBFFFC00000016FFDBBFFB965A5B3FA1F5E0FFC00001;
defparam sdpb_inst_2.INIT_RAM_2E = 256'hFC7DFF9E56FE41053FFE19772621FF7DD60000004749D51FFF1EDF7BD7FFEFB8;
defparam sdpb_inst_2.INIT_RAM_2F = 256'hFFFFA13125DFFFE6DFFFC80A3FFFE39C633E7128F10000000600407FFFE430D9;
defparam sdpb_inst_2.INIT_RAM_30 = 256'h0000E979FFFFFF9CBCF7EFFDADFFC200EDFFFE1C07705880FA000000010018D5;
defparam sdpb_inst_2.INIT_RAM_31 = 256'h314E000000F7EE01FFFFFFF3BBDE7BF6F2BFFD0046FFFFD0FF19E7A0DD800000;
defparam sdpb_inst_2.INIT_RAM_32 = 256'hF869883E08036000B780603FFFFFFFFF87FFFF7FFB5FFF2043DFBEFF018528F0;
defparam sdpb_inst_2.INIT_RAM_33 = 256'h26EEF1F7FE12335E0206100166A00003FFFDFFFFE4377DDFFFF5FF941F2F557F;
defparam sdpb_inst_2.INIT_RAM_34 = 256'h77DEFFFE055AE63BF78D2937D1A7F30268E000000242D3FFFEE7CB3FFDF7BFF1;
defparam sdpb_inst_2.INIT_RAM_35 = 256'hFFFB1D56FF7FE7FFE1445EE37FF292FDE3D0FAE7AEC0005F508B267FFFDE7BFF;
defparam sdpb_inst_2.INIT_RAM_36 = 256'hE0344697FFFF43EADFFEC7FFE07E20C987F88B82FC4C7F7FBBC48E22E0510F7F;
defparam sdpb_inst_2.INIT_RAM_37 = 256'hD9F2742E80146A107FFFF38D6BFFE7FFFA1C9338EFFC5B197EA61FDFA5CC199C;
defparam sdpb_inst_2.INIT_RAM_38 = 256'h47F9B2EB09FEE7CE00063D4B33DBFEFDA47FFFFFFE4B6032011F98059F90C0CB;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h4003F53E23F2672117DFEB7A0004D4014C3BFFD6431FE77FFE407F5A005FCAEA;
defparam sdpb_inst_2.INIT_RAM_3A = 256'hFDE20161C025F93D93FF27A5B4FBEBBC000103FFF483FFFBC253FFDEF7A81D40;
defparam sdpb_inst_2.INIT_RAM_3B = 256'hEB04F7FDFFF900980807FCCBB9F7BBFDFD7EF4E8800058FFFF79EFFF1A5EBFEF;
defparam sdpb_inst_2.INIT_RAM_3C = 256'hFFFF6DFFFC5F20FF73BF93B20009FC5D2C3FFBFFEFBFEB7F40006A3FFFF3BFFF;
defparam sdpb_inst_2.INIT_RAM_3D = 256'hCC000AE37FFFE9FFFF95EDDFFFFF808E9EDBFF27013FFFBFEC1FE67FC4001F9F;
defparam sdpb_inst_2.INIT_RAM_3E = 256'hFE87F27FFE4002F03FFFFABFFFC2E7E3FFFBDA297CA03F92EA9FFEFFFB07F37F;
defparam sdpb_inst_2.INIT_RAM_3F = 256'h8813FFFFFEDBF93FFFEC43EC0FFFFE3FFFF443E57FFF7B02DFFFFBCEF7A3FF7F;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[3]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b1;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'hFFFFFFE08066FDFBFFFFFFFE800000000FFFFFFFFFFEDCFE5FFFFFFFFFFFFE42;
defparam sdpb_inst_3.INIT_RAM_01 = 256'h10777FFFFFFFFFFC0003B3FFFFFFFFFE000280001C7FFFFFFEFBF7FF5BFFFFFF;
defparam sdpb_inst_3.INIT_RAM_02 = 256'hE90000042BDC377FFFFFFFFF441BFFFFFFFFFFFE0005F000006CEEDBFF460058;
defparam sdpb_inst_3.INIT_RAM_03 = 256'h00013BE42C000800082523FFFFFFFFFFB803FEFFFFFFFFFF4003FE00000DAF85;
defparam sdpb_inst_3.INIT_RAM_04 = 256'h0001FFE2800101B082100000000301FFFFFFFFFFFF0FFFFFFFFFFFFF0000FFC0;
defparam sdpb_inst_3.INIT_RAM_05 = 256'hFFFFFFFF8081E5FFF80245BE28300000007871F9FFFFFFFFFFA3FFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_06 = 256'hFFFFFF7FFFFFFFFFFE03FF59FF8070DFF4400210000221AFFFFFFFFFFFFDFFFF;
defparam sdpb_inst_3.INIT_RAM_07 = 256'hF7FFFFFFFFFFFFFFFFFFFFFFFE00FFEFFFFFF6B7FEC30080020000167FFFFFFF;
defparam sdpb_inst_3.INIT_RAM_08 = 256'h0840001EFFFFFFFFFFFFFFFDBFFFFFFFFF10FFFD7FF7FFFFFF6000505000100D;
defparam sdpb_inst_3.INIT_RAM_09 = 256'hFFFE0000C0800005397FFFFFFFFFFDFFFFFFFFFFFFC81BFB7DEFFFFFFFFC0008;
defparam sdpb_inst_3.INIT_RAM_0A = 256'hFFFEFFEFFFFB0007A74018100FDFFFFFFFFFFF7FFFFFFFFFFFE81FFEFFE9FF7F;
defparam sdpb_inst_3.INIT_RAM_0B = 256'hFFFF7FFFBFF42FD3FFFE820302E0000013FDFFFFFFFFFFBFFDFFFFFFFFFFFFDA;
defparam sdpb_inst_3.INIT_RAM_0C = 256'hFFFFFFFFFFFFCFFC29FA6AEBFFFFC0039214000000FEFFFFEFDFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0D = 256'hBFFFFFFFFFFFFFFFFFFFF8FE7D79FF29FFFFF400C54E2000007F1DF6FFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_0E = 256'h0001E39DFE73FFFFFFFFFFFFFFFFFE8E1F8F7FE1FFFFF9006961FC00004AFFFE;
defparam sdpb_inst_3.INIT_RAM_0F = 256'h0F58027200800DF6F6DFFFFFFFFFFFFFFFFFFFFC3FF3CFF9FDFFFF0019109B00;
defparam sdpb_inst_3.INIT_RAM_10 = 256'hFFA1FFF801EC07EE0064002BBF5FFBFFFFFFFFFFFFFFFFF78FFC197EBFFFFFC0;
defparam sdpb_inst_3.INIT_RAM_11 = 256'hFDBFCFD977B03FF340BF0CAFC0001012FEBF7FFFFFFBFFFFFFFFFFFDE3FE8DBD;
defparam sdpb_inst_3.INIT_RAM_12 = 256'hFFFFFFFFEFB307FD9FE607FF602F405F7400801D5FFEF1FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_13 = 256'hC6FFFFFFFFFFFFFFFECFEDFEABD7C0FFFBFFE1FCFF0000103FBCD6C1B1FFFFFF;
defparam sdpb_inst_3.INIT_RAM_14 = 256'h50F6F1D7BD1FFFFFFFFFFFFFFF69FAF773EBDC3FFFFFFD5DE7E00001CA6BBA77;
defparam sdpb_inst_3.INIT_RAM_15 = 256'h15F1800002FFFFA337FFFFFFFFFFFFFFFFD93EBF85F1F70FFFFDFF96E75C0000;
defparam sdpb_inst_3.INIT_RAM_16 = 256'hFFE3B37763AF3800004BEFFEBFBFFF7FFFFFFFFFFFFF0F68C3593FE3FFF54FF3;
defparam sdpb_inst_3.INIT_RAM_17 = 256'h35ECFF663FE7DD324D7C674000077EDFD9FFFFFFFFFFFFFFFFFDFFDFBDE6DE39;
defparam sdpb_inst_3.INIT_RAM_18 = 256'hF7FFCDFB43FCFEA907E7B398CDE2E7F00001FFF9A43BFFFFFFFFFFFFFFFFBCBC;
defparam sdpb_inst_3.INIT_RAM_19 = 256'hFFFFFFE7FE7FE363C89F9F9A83F3B9F90524BB7F0006FFFFE43FFDFFFFFFFFFF;
defparam sdpb_inst_3.INIT_RAM_1A = 256'hFFF3B5BFFFFFFFFFBA3B78F3FC27979C80FCE70045441FD3F50877FF3A1535FF;
defparam sdpb_inst_3.INIT_RAM_1B = 256'h745553FFFFD113DFFFFFFFFF0F0E9E167C7DFDEF107E2FBFE79C05DF3F4007FF;
defparam sdpb_inst_3.INIT_RAM_1C = 256'hFFE1C29FA3F99FD7FE61AB5FDFFFFFF6C1F7D30227F4AE5DE60F3CCFFE0A00CD;
defparam sdpb_inst_3.INIT_RAM_1D = 256'hFA700141FFF8415BC6C07FFFF956557BE7FFFFFFBA58FBC002FE4FFF54C30E77;
defparam sdpb_inst_3.INIT_RAM_1E = 256'hEE0C74F3F91C008C7FFF50620BD786FFFDC6545E7BFFFFFF811E3DE1C03BE7F5;
defparam sdpb_inst_3.INIT_RAM_1F = 256'hFFC00FF87339BF3E780E00289FFFD95D1F87FCFFFFFFDFC9BFFFFFFFFCC33630;
defparam sdpb_inst_3.INIT_RAM_20 = 256'h8FEFFFFFFFF00FF83C64F4EFC9C3810E17FFF6E7B36FFF97FEFF86C9BFFBFFFF;
defparam sdpb_inst_3.INIT_RAM_21 = 256'hFFF7F6E7BAF8FFFFFFFE03AF1E1FFDF6FAE1C001A4FFFA01E827FFD2FFFFE07C;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h1E993FFBD7FFC494B11E7FFFFF7F47138F03FE7FBCF8E03E6F9FFC657A43FFFE;
defparam sdpb_inst_3.INIT_RAM_23 = 256'hD0547E3CDF81EFFFC4FFEFCE427F8F7FFFBFFCD80700610D5F1878018937FE35;
defparam sdpb_inst_3.INIT_RAM_24 = 256'h17BE1F00BE7E8156E7E43FFFF9BFFDBFE579E3FFFFED9076488000076F0C1E01;
defparam sdpb_inst_3.INIT_RAM_25 = 256'h79D8E07E1BCE1F003F82FF561BFDB7BFF0C7FFFCB4FEF8EFFFD9200F230F8000;
defparam sdpb_inst_3.INIT_RAM_26 = 256'hFFECA002F106187FF1B01FC04FF2BEEC13FF40FBF075FFF9F5B99E7FFBFFC00F;
defparam sdpb_inst_3.INIT_RAM_27 = 256'hDDC03FE3FFF7E800C201B63FFFB5FFC03FFE49A6B9FFC9C3803F7FF5F7BBBF83;
defparam sdpb_inst_3.INIT_RAM_28 = 256'hF348A7FFF8D027F9FFFFCE0020C0B59FFEF03EC00FFFE4A941FFFAFD3FFCDFF7;
defparam sdpb_inst_3.INIT_RAM_29 = 256'h7DFFFFCB15E4BDFFFC3101FE3FFFEC801E30A567D100000003FFFC5673FFFE5E;
defparam sdpb_inst_3.INIT_RAM_2A = 256'h01FFFFFFE0FFB3F9108CBF7FFFF2B0C79FFFFFC007008513E000000002FFFFE0;
defparam sdpb_inst_3.INIT_RAM_2B = 256'h7000000005FFFFFFFFFFFFFF149EFECFFEF3C38FE4BFFBC001CAF1A8E0000000;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h401F21C93800000008FFFFFFFFFFFF7FF3A5BEFBFEF677F8F8FFFFD6007B8736;
defparam sdpb_inst_3.INIT_RAM_2D = 256'hFF8DFFFCC000E7D31E00040003FFFFFFFFFFFFBFFC18C37FFFA1F5E0FE3FFFFE;
defparam sdpb_inst_3.INIT_RAM_2E = 256'hADFDFF9E56E1BEFAC0001E7F1E20008229FFFFFFFFFFE7FFFFE0E67FFFFFEFB8;
defparam sdpb_inst_3.INIT_RAM_2F = 256'hFFFFFE757FBFFFE6DFF837F5C00003E01F3E0ED70EFFFFFFFFFFF3E7FFFFC3FB;
defparam sdpb_inst_3.INIT_RAM_30 = 256'hFFFE3D07FFFFFFECBCEFEFFDADFE3DFF1200001FFFCFC77F05FFFFFFFFFFCBD3;
defparam sdpb_inst_3.INIT_RAM_31 = 256'hC7E1FFFFFF32E9FFFFFFFFFD9ADEFBF6F2BF82FFB9000000FFEE105F227FFFFF;
defparam sdpb_inst_3.INIT_RAM_32 = 256'h0076AB01F7FD1FFF4AE61FFFFFFFFFFFC3FF9F7FFB5FE0DFBC20410001F28C0F;
defparam sdpb_inst_3.INIT_RAM_33 = 256'hD9110E080019C041FDF9F7FE8B1FFFFFFFFFFFFFF8BF3FDFFFF5F86BE0D0AA00;
defparam sdpb_inst_3.INIT_RAM_34 = 256'h77DEFF81FAA519C4080F29D02ED80CFDBB1FFFFFFFFCB3FFFF37DD7FFDF7BE0E;
defparam sdpb_inst_3.INIT_RAM_35 = 256'hFFFC596DFF7FE7E01EBBA11C8003658C1C3F0518343FFF8CAF7FFAFFFFE6FFEF;
defparam sdpb_inst_3.INIT_RAM_36 = 256'h1FC0D1FFFFFFABF73FFEC7F81F81DF367800F24603BF80E0523B708D5F9E5DBF;
defparam sdpb_inst_3.INIT_RAM_37 = 256'h640D87A17FE5DAD07FFFFEC737FFE7FE05E36CC7100068730159E0200033E244;
defparam sdpb_inst_3.INIT_RAM_38 = 256'hC0064D1C74010001FFFE12FB03DBFFDFDBFFFFFF81B49FCDFEE01581806F3F38;
defparam sdpb_inst_3.INIT_RAM_39 = 256'hBFFC0636600D9BD802200845FFF813FE407BFFFBF8DFE77FE1BF80A5FFA00C70;
defparam sdpb_inst_3.INIT_RAM_3A = 256'hFE1DFE9E3FDA014AB000D83C06040203FFFE07FFF987FFFF7E8FFFDEF857E2BF;
defparam sdpb_inst_3.INIT_RAM_3B = 256'hFDCD0FFDFF86FF67F7F800BBE808440C390119977FFF6FFFFFAA6FFFAD80FFEF;
defparam sdpb_inst_3.INIT_RAM_3C = 256'hFFFFCBFFFEA0DFFF73E06C4DFFF60077B40004000C800200BFFF83FFFFF92FFF;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h33FFF01FFFFFFC3FFFC0927FFFF87F7161240036D30000400B8003003BFFEC7F;
defparam sdpb_inst_3.INIT_RAM_3E = 256'h03A0000001BFFC67FFFFFC8FFFF8170FFFFE25D6835FC01ABF80010001C00900;
defparam sdpb_inst_3.INIT_RAM_3F = 256'h7330000000A800000013BC67FFFFFFA9FFFF522AFFFF84FD2000040F4A600080;

SDPB sdpb_inst_4 (
    .DO({sdpb_inst_4_dout_w[30:0],sdpb_inst_4_dout[4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[4]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_4.READ_MODE = 1'b1;
defparam sdpb_inst_4.BIT_WIDTH_0 = 1;
defparam sdpb_inst_4.BIT_WIDTH_1 = 1;
defparam sdpb_inst_4.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_4.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_4.RESET_MODE = "SYNC";
defparam sdpb_inst_4.INIT_RAM_00 = 256'hFFFFFFFF7FFFFFFFFFFFFFFE800000000FFFFFFFFFFEDCFE5FFFFFFFFFFFFFFC;
defparam sdpb_inst_4.INIT_RAM_01 = 256'h10777FFFFFFFFFFFFFFFFFFFFFFFFFFE000080001C7FFFFFFEFBF7FF5BFFFFFF;
defparam sdpb_inst_4.INIT_RAM_02 = 256'hE90000042BDC377FFFFFFFFFFFFFFFFFFFFFFFFE0007F000006CEEDBFF460058;
defparam sdpb_inst_4.INIT_RAM_03 = 256'h00013BE42C000800082523FFFFFFFFFFFFFFFFFFFFFFFFFF4003FF00000DAF85;
defparam sdpb_inst_4.INIT_RAM_04 = 256'h00015FFB800101B082100000000301FFFFFFFFFFFFFFFFFFFFFFFFFF0001FFF0;
defparam sdpb_inst_4.INIT_RAM_05 = 256'hFFFFFFFF80816FE9F80245BE28300000007871F9FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFE037FEDFF8070DFF4400210000221AFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_07 = 256'hF7FFFFFFFFFFFFFFFFFFFFFFFE00FFE4FFDFF6B7FEC30080020000167FFFFFFF;
defparam sdpb_inst_4.INIT_RAM_08 = 256'h0840001EFFFFFFFFFFFFFFFFFFFFFFFFFF10BFF77FFBFFFFFF6000505000100D;
defparam sdpb_inst_4.INIT_RAM_09 = 256'hFFFE0000C0800005397FFFFFFFFFFFFFFFFFFFFFFFC84BFEF7EBFFFFFFFC0008;
defparam sdpb_inst_4.INIT_RAM_0A = 256'h7FF4FFD7FFFB0007EB4018100FDFFFFFFFFFFFFFFFFFFFFFFFE81CBFFF7FFF7F;
defparam sdpb_inst_4.INIT_RAM_0B = 256'hFFFF7FFE7FF76FDDFFFE8203AFE0000013FDFFFFFFFFFFFFFFFFFFFFFFFFDFEB;
defparam sdpb_inst_4.INIT_RAM_0C = 256'hFFFFFFFFFFFFDFFD99FB77F97FFFC003635C000000FEFFFFEFDFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0D = 256'hBFFFFFFFFFFFFFFFFFFFFBFF9E7B7EEFDFFFF400B742A000007F1DF6FFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_0E = 256'h0001E39DFE73FFFFFFFFFFFFFFFFFF3EDFBDFFEEF7FFF9006F79EC00004AFFFE;
defparam sdpb_inst_4.INIT_RAM_0F = 256'h0FE3FFF200800DF6F6DFFFFFFFFFFFFFFFFFFFF75FF28FFF7DFFFF001FA3FF00;
defparam sdpb_inst_4.INIT_RAM_10 = 256'h77BFFFF801FFFBCE0064002BBF5FFBFFFFFFFFFFFFFFFFF72FFDE97D1F7FFFC0;
defparam sdpb_inst_4.INIT_RAM_11 = 256'hFFEF6FE8FD9FFFF340BDFC01C0001012FEBF7FFFFFFFFFFFFFFFFFFDEFFE4EBD;
defparam sdpb_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFB627FEFF3DFFFF602F88003400801D5FFEF1FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_13 = 256'hC6FFFFFFFFFFFFFFFECF75FEDFCF3FFFFBFFF0910F0000103FBCD6C1B1FFFFFF;
defparam sdpb_inst_4.INIT_RAM_14 = 256'h50F6F1D7BD1FFFFFFFFFFFFFFF3FF2F70FE7C3FFFFFFFE1128E00001CA6BBA77;
defparam sdpb_inst_4.INIT_RAM_15 = 256'h801F800002FFFFA337FFFFFFFFFFFFFFFFDE7FEFA4F4F0FFFFFEFFEA063C0000;
defparam sdpb_inst_4.INIT_RAM_16 = 256'hFFF28DBFB100F800004BEFFEBFBFFFFFFFFFFFFFFFFF7FFEFF1B7C1FFFFD67FD;
defparam sdpb_inst_4.INIT_RAM_17 = 256'hF1FF72E1FFFCB06E76239F4000077EDFD9FFFFFFFFFFFFFFFFFFF7DFF3E4CC87;
defparam sdpb_inst_4.INIT_RAM_18 = 256'hEFFFFBBFFF7DFCE8FFFBF42F6ECD40F00001FFF9A43BFFFFFFFFFFFFFFFFFEFD;
defparam sdpb_inst_4.INIT_RAM_19 = 256'hFFFFFFF5FF7FFDF7AFBE7FDA7FFD64037AC1603F0006FFFFE43FFDFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_1A = 256'hFFF3B5BFFFFFFFFBFFFFFF69F9EFFFAC7FFFF6FF9BF8A103F50877FF3A1535FF;
defparam sdpb_inst_4.INIT_RAM_1B = 256'h867553FFFFD113DFFFFFFFFFF7FEFFFFFF9B9BF34FFF9D7FFAEB90107F4007FF;
defparam sdpb_inst_4.INIT_RAM_1C = 256'hFFF5FC410BFB9FD7FE61AB5FFFFFFFFFFFFFABFFDF318FCCE1FFD63FFF9CF210;
defparam sdpb_inst_4.INIT_RAM_1D = 256'hCA0FFCA7FFFE7B880FBFEFFFF956557BFFFFFFFFDDBF6FFF7AFF3FD7843FF52F;
defparam sdpb_inst_4.INIT_RAM_1E = 256'h0E9E7DF3F903FF1DFFFFAFF90FDFFFFFFDC6545E7FFFFFFF7FA0CBFE1ECBF3E1;
defparam sdpb_inst_4.INIT_RAM_1F = 256'hFFFFF00F83FFBF787C01FFD7FFFFEBFE3FFFFFFFFFFFDFC9BFFFFFFFF33CC9FF;
defparam sdpb_inst_4.INIT_RAM_20 = 256'h8FFFFFFFFFF7F003C07DF1DEC9C07FF5EFFFFBBFD7FFFFF3FEFF86C9BFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_21 = 256'hFFF7F6E7BAFFFFFFFFFFFC2FE01FFEECF9E03FFE1FFFFC7BF3FFFFFFFFFFE07C;
defparam sdpb_inst_4.INIT_RAM_22 = 256'h7F3FFFFFDFFFC494B11FFFFFFFFFFC607003FEFFFFF81FFFBBFFFF08FCDBFFFF;
defparam sdpb_inst_4.INIT_RAM_23 = 256'hFE0BFFF17FEDFFFFFFFFEFCE427FFFFFFFFFFFE5FC00611FFF9807FFF56FFFBA;
defparam sdpb_inst_4.INIT_RAM_24 = 256'h1E9E00FFFFA0FEA5FFFB3FFFFFFFFDBFE579FFFFFFFFFFFFFF000003EF0C01FF;
defparam sdpb_inst_4.INIT_RAM_25 = 256'h09F3E000199E00FFFFF7DDF9B7FEAFFFFFDFFFFCB4FEFFFFFFFFFFFF23FF8000;
defparam sdpb_inst_4.INIT_RAM_26 = 256'hFFFFFFFDE3FCF8000180003FFFFCA57217FF9DFFFFF3FFF9F5B99FFFFFFFFFF7;
defparam sdpb_inst_4.INIT_RAM_27 = 256'hDDC03FFFFFFFFFFF57FF0E00000E003FFFFF81DDD7FFF27EFFFAFFF5F7BBBFFF;
defparam sdpb_inst_4.INIT_RAM_28 = 256'hEF77FFFFF8D027FFFFFFFFFFC87FD380010FC13FFFFFF953EFFFFC87FFFEBFF7;
defparam sdpb_inst_4.INIT_RAM_29 = 256'h83FFFFF2DFFB03FFFC3101FFFFFFFFFFE13FACE02EFFFFFFFFFFFF9FAFFFFF90;
defparam sdpb_inst_4.INIT_RAM_2A = 256'hFFFFFFFFFFFFB3FE348B80FFFFF2B0C7FFFFFFFFF8237F701FFFFFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2B = 256'h0FFFFFFFFFFFFFFFFFFFFFFFE6DD003FFEF3C38FFFFFFFFFFE0EFD181FFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2C = 256'hFFE0338707FFFFFFFFFFFFFFFFFFFF7FFC384087FEF677F8FFFFFFFFFF83D8EE;
defparam sdpb_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFF064F01FFFFFFFFFFFFFFFFFFFFBFFFE08484FFA1F5E0FFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_2E = 256'h51FDFF9E56FFFFFFFFFFE07F01DFFFFFFFFFFFFFFFFFFAFFFFFF0A863FFFEFB8;
defparam sdpb_inst_4.INIT_RAM_2F = 256'hFFFFFFA2D03FFFE6DFFFFFFFFFFFFC0000C1FFFFFFFFFFFFFFFFFBEFFFFFFD4C;
defparam sdpb_inst_4.INIT_RAM_30 = 256'hFFFFC0FFFFFFFFF64007EFFDADFFFFFFFFFFFFE000303FFFFFFFFFFFFFFFE54F;
defparam sdpb_inst_4.INIT_RAM_31 = 256'hFBDFFFFFFFC0C7FFFFFFFFFEC129FBF6F2BFFFFFFFFFFFFF000F0FFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_32 = 256'hFF879AFFFBFFFFFFFC11FFFFFFFFFFFFE8003F7FFB5FFFFFFFFFFFFFFE1F9BFF;
defparam sdpb_inst_4.INIT_RAM_33 = 256'hFFFFFFFFFFE1843FFFFFFFFFF97FFFFFFFFFFFFFFD4027DFFFF5FFFFFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_34 = 256'h77DEFFFFFFFFFFFFFFF1E2CFFF7FFFFFD0FFFFFFFFFF17FFFF88A47FFDF7BFFF;
defparam sdpb_inst_4.INIT_RAM_35 = 256'hFFFEA401FF7FE7FFFFFFFFFFFFFC3F63FFDFFF7FE9FFFFF3FFFFFFFFFFF1040F;
defparam sdpb_inst_4.INIT_RAM_36 = 256'hFFFCD3FFFFFFD4083FFEC7FFFFFFFFFFFFFF3DB1FFF7FFDF91FFFF36C01DEB7F;
defparam sdpb_inst_4.INIT_RAM_37 = 256'hCBFFFB5FFFF5FED07FFFF800C7FFE7FFFFFFFFFFFFFF88F8FFFEFFFFCBFFFCD3;
defparam sdpb_inst_4.INIT_RAM_38 = 256'h3FFFF7FB8BFFFA3FFFFA30FF83DBFF0104FFFFFFFFFFFFFFFFFFE4047FFFBFFF;
defparam sdpb_inst_4.INIT_RAM_39 = 256'hFFFFF82F1FFFFDFBD9FFF63FFFFE0FFF847BFFE04A1FE77FFFFFFFFFFFFFF2F2;
defparam sdpb_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFE4F0FFFFFFBEDFFF67FFFFF0FFFFF87FFFC0927FFDEFFFFFFFF;
defparam sdpb_inst_4.INIT_RAM_3B = 256'hF0350FFDFFFFFFFFFFFFFF3D27FFFFF7CCFFE77FFFFFCBFFFFD86FFFC0307FEF;
defparam sdpb_inst_4.INIT_RAM_3C = 256'hFFFFABFFFF0047FF73FFFFFFFFFFFF97B3FFFFFFF27FFCFFFFFFC1FFFFFF8FFF;
defparam sdpb_inst_4.INIT_RAM_3D = 256'hFFFFFC3FFFFFF47FFFE0043FFFFFFFFFFFFFFFCB78FFFFFFF37FFEFFFFFFF4FF;
defparam sdpb_inst_4.INIT_RAM_3E = 256'hFC5FFAFFFFFFFF6FFFFFFE9FFFFC0107FFFFFFFFFFFFFFE3A27FFFFFFFBFF4FF;
defparam sdpb_inst_4.INIT_RAM_3F = 256'hEF8FFFFFFF07FF7FFFFFFFA7FFFFFFF9FFFF8228FFFFFFFFFFFFFFF3DB1FFFFF;

SDPB sdpb_inst_5 (
    .DO({sdpb_inst_5_dout_w[30:0],sdpb_inst_5_dout[5]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_5.READ_MODE = 1'b1;
defparam sdpb_inst_5.BIT_WIDTH_0 = 1;
defparam sdpb_inst_5.BIT_WIDTH_1 = 1;
defparam sdpb_inst_5.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_5.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_5.RESET_MODE = "SYNC";
defparam sdpb_inst_5.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFE800000000FFFFFFFFFFEDCFE5FFFFFFFFFFFFFFE;
defparam sdpb_inst_5.INIT_RAM_01 = 256'h10777FFFFFFFFFFFFFFFFFFFFFFFFFFE000080001C7FFFFFFEFBF7FF5BFFFFFF;
defparam sdpb_inst_5.INIT_RAM_02 = 256'hE90000042BDC377FFFFFFFFFFFFFFFFFFFFFFFFE00061000006CEEDBFF460058;
defparam sdpb_inst_5.INIT_RAM_03 = 256'h00013BE42C000800082523FFFFFFFFFFFFFFFFFFFFFFFFFF40020100000DAF85;
defparam sdpb_inst_5.INIT_RAM_04 = 256'h0001E01C800101B082100000000301FFFFFFFFFFFFFFFFFFFFFFFFFF00000030;
defparam sdpb_inst_5.INIT_RAM_05 = 256'hFFFFFFFF80819E0E080245BE28300000007871F9FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFE0380FE008070DFF4400210000221AFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_07 = 256'hF7FFFFFFFFFFFFFFFFFFFFFFFE00801F001FF6B7FEC30080020000167FFFFFFF;
defparam sdpb_inst_5.INIT_RAM_08 = 256'h0840001EFFFFFFFFFFFFFFFFFFFFFFFFFF10C00EE018FFFFFF6000505000100D;
defparam sdpb_inst_5.INIT_RAM_09 = 256'hFFFE0000C0800005397FFFFFFFFFFFFFFFFFFFFFFFC87C078E0C0FFFFFFC0008;
defparam sdpb_inst_5.INIT_RAM_0A = 256'h800F001FFFFB0007D74018100FDFFFFFFFFFFFFFFFFFFFFFFFE823C700EC007F;
defparam sdpb_inst_5.INIT_RAM_0B = 256'hFFFF6003C00EE03FFFFE82039360000013FDFFFFFFFFFFFFFFFFFFFFFFFFE03F;
defparam sdpb_inst_5.INIT_RAM_0C = 256'hFFFFFFFFFFFFD003FE031F0EFFFFC003834C000000FEFFFFEFDFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0D = 256'hBFFFFFFFFFFFFFFFFFFFFF00C30781EC3FFFF400C321A000007F1DF6FFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_0E = 256'h0001E39DFE73FFFFFFFFFFFFFFFFFF71E079801E0FFFF90072AA1C00004AFFFE;
defparam sdpb_inst_5.INIT_RAM_0F = 256'h0F94017200800DF6F6DFFFFFFFFFFFFFFFFFFFF3E00FF00603FFFF001C040300;
defparam sdpb_inst_5.INIT_RAM_10 = 256'hC01FFFF801F607DE0064002BBF5FFBFFFFFFFFFFFFFFFFF77003DE83407FFFC0;
defparam sdpb_inst_5.INIT_RAM_11 = 256'hFC70F03E805FFFF340BE8481C0001012FEBF7FFFFFFFFFFFFFFFFFFFE701F3C3;
defparam sdpb_inst_5.INIT_RAM_12 = 256'hFFFFFFFFFFBFF803C04BFFFF602FD4187400801D5FFEF1FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_13 = 256'hC6FFFFFFFFFFFFFFFCCFFA01C000FFFFFBFFFB90070000103FBCD6C1B1FFFFFF;
defparam sdpb_inst_5.INIT_RAM_14 = 256'h50F6F1D7BD1FFFFFFFFFFFFFFF19FF08F8103FFFFFFFFFB108E00001CA6BBA77;
defparam sdpb_inst_5.INIT_RAM_15 = 256'h821B800002FFFFA337FFFFFFFFFFFFFFFFF87C7078010FFFFFFF3FF6171C0000;
defparam sdpb_inst_5.INIT_RAM_16 = 256'hFFF440AFD1107800004BEFFEBFBFFFFFFFFFFFFFFFFF5FB710A041FFFFFEB1FE;
defparam sdpb_inst_5.INIT_RAM_17 = 256'hFC0404BFFFF907853A210F4000077EDFD9FFFFFFFFFFFFFFFFFEF1CF780402FF;
defparam sdpb_inst_5.INIT_RAM_18 = 256'hFFFFF7B87E8300DFFFFC0C2C374161F00001FFF9A43BFFFFFFFFFFFFFFFFFED9;
defparam sdpb_inst_5.INIT_RAM_19 = 256'hFFFFFFF5FF7FFF27CFC140A7FFFE1BFD62F0011F0006FFFFE43FFDFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_1A = 256'hFFF3B5BFFFFFFFFFFFDFFFE1F7F030037FFF0DFFECBE0103F50877FF3A1535FF;
defparam sdpb_inst_5.INIT_RAM_1B = 256'h8CB553FFFFD113DFFFFFFFFEFFF7FFFE3D580030BFFFC2FFFC07C020FF4007FF;
defparam sdpb_inst_5.INIT_RAM_1C = 256'hFFFA1F0304049FD7FE61AB5FFFFFFFF7DFFBFBFBC73E51283FFFE97FFFD37812;
defparam sdpb_inst_5.INIT_RAM_1D = 256'h25FFFE0FFFFF47E000409FFFF956557BFFFFFFFFFFFF7DFF736FC040ABFFF9DF;
defparam sdpb_inst_5.INIT_RAM_1E = 256'hF0BF7F0A06FFFF83FFFFC1FC08A001FFFDC6545E7FFFFFFF7DB8FBFFEED7EC1A;
defparam sdpb_inst_5.INIT_RAM_1F = 256'hFFFFFFEFFC1F8F8147FFFFE87FFFF43F9000001FFFFFDFC9BFFFFFFFFFFFFFBF;
defparam sdpb_inst_5.INIT_RAM_20 = 256'h8FFFFFFFFFFFFFFBFF83FAC2043FFFFA1FFFFD4FE200000FFEFF86C9BFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_21 = 256'h3FF7F6E7BAFFFFFFFFFFFFD17FE00CD2821FFFFF47FFFF87FD800000FFFFE07C;
defparam sdpb_inst_5.INIT_RAM_22 = 256'hFFD8000027FFC494B11FFFFFFFFFFFFC0FFC003C0307FFFFD07FFFD5FF440000;
defparam sdpb_inst_5.INIT_RAM_23 = 256'hFF63FF96BFF4000001FFEFCE427FFFFFFFFFFF3E03FF9EEFC0E7FFFFFADFFFE1;
defparam sdpb_inst_5.INIT_RAM_24 = 256'hDD41FFFFFFDB7F881FFD4000007FFDBFE579FFFFFFFFFF80007FFFFDE0B3FFFF;
defparam sdpb_inst_5.INIT_RAM_25 = 256'hF60C1FFFE741FFFFFFF80680AFFF1000003FFFFCB4FEFFFFFFFFFFC0DC207FFF;
defparam sdpb_inst_5.INIT_RAM_26 = 256'hFFFFFFFF1C0207FFFE4FFFFFFFFFC2018FFFEA00000FFFF9F5B99FFFFFFFFFF0;
defparam sdpb_inst_5.INIT_RAM_27 = 256'hDDC03FFFFFFFFFFFAC0081FFFFFFFFFFFFFFEE044FFFFD010007FFF5F7BBBFFF;
defparam sdpb_inst_5.INIT_RAM_28 = 256'h00801FFFF8D027FFFFFFFFFFFF80707FFFFFFFFFFFFFFEE4DFFFFF2800037FF7;
defparam sdpb_inst_5.INIT_RAM_29 = 256'hFFFFFFFCA00087FFFC3101FFFFFFFFFFFDC06C1FFFFFFFFFFFFFFFE01FFFFFE5;
defparam sdpb_inst_5.INIT_RAM_2A = 256'hFFFFFFFFFFFFB3FFD97080FFFFF2B0C7FFFFFFFFFFCEFB0FFFFFFFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF8E8001FFEF3C38FFFFFFFFFFFF3F887FFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2C = 256'hFFFFC3E0FFFFFFFFFFFFFFFFFFFFFF7FFFC08003FEF677F8FFFFFFFFFFFC3721;
defparam sdpb_inst_5.INIT_RAM_2D = 256'hFFFFFFFFFFFFF8C0FFFFFFFFFFFFFFFFFFFFFFBFFFFF20007FA1F5E0FFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_2E = 256'h53FDFF9E56FFFFFFFFFFFF80FFFFFFFFFFFFFFFFFFFFFC3FFFFFF6002FFFEFB8;
defparam sdpb_inst_5.INIT_RAM_2F = 256'hFFFFFFD0027FFFE6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF81FFFFFFEC0;
defparam sdpb_inst_5.INIT_RAM_30 = 256'hFFFF0BFFFFFFFFFA030FEFFDADFFFFFFFFFFFFFFFF87FFFFFFFFFFFFFFFFF37F;
defparam sdpb_inst_5.INIT_RAM_31 = 256'hFFCFFFFFFFE85FFFFFFFFFFF4001FBF6F2BFFFFFFFFFFFFFFFF27FFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_32 = 256'hFFFAA1FFFFFFFFFFFE2FFFFFFFFFFFFFF8043F7FFB5FFFFFFFFFFFFFFFFCE7FF;
defparam sdpb_inst_5.INIT_RAM_33 = 256'hFFFFFFFFFFFF56FFFFFFFFFFF9FFFFFFFFFFFFFFFF1027DFFFF5FFFFFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_34 = 256'h77DEFFFFFFFFFFFFFFFEC8BFFFFFFDFFE5FFFFFFFFFFC7FFFFE0047FFDF7BFFF;
defparam sdpb_inst_5.INIT_RAM_35 = 256'hFFFF8611FF7FE7FFFFFFFFFFFFFF865FFFFFFFFFCBFFFFFA000001FFFFFC020F;
defparam sdpb_inst_5.INIT_RAM_36 = 256'hFFFB2C07FFFFF0083FFEC7FFFFFFFFFFFFFFCE2FFFFFFFFFC7FFFF4A3FE008FF;
defparam sdpb_inst_5.INIT_RAM_37 = 256'h87FFFCBFFFFA012FBFFFFE10C7FFE7FFFFFFFFFFFFFFF717FFFEFFEF87FFFF0F;
defparam sdpb_inst_5.INIT_RAM_38 = 256'hFFFFF7FFC7FFFD7FFFFDCF007DDBFFC104FFFFFFFFFFFFFFFFFFFBF3FFFFFFF7;
defparam sdpb_inst_5.INIT_RAM_39 = 256'hFFFFFEF2FFFFFFFFD7FFF9FFFFFFFFFFFBFBFFF94A1FE77FFFFFFFFFFFFFFD29;
defparam sdpb_inst_5.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFB37FFFFFBBC3FFF8FFFFFFFFFFFE7FFFFF0C27FFDEFFFFFFFF;
defparam sdpb_inst_5.INIT_RAM_3B = 256'hFC159FFDFFFFFFFFFFFFFFC69FFFFFFBEBFFF0FFFFFFB7FFFFE7EFFFE410FFEF;
defparam sdpb_inst_5.INIT_RAM_3C = 256'hFFFFD7FFFF8045FF73FFFFFFFFFFFFE96FFFFFFFF1FFFBFFFFFFFFFFFFFC7FFF;
defparam sdpb_inst_5.INIT_RAM_3D = 256'hFFFFFFFFFFFFFBFFFFF0063FFFFFFFFFFFFFFFF497FFFFFFFEFFF3FFFFFFFBFF;
defparam sdpb_inst_5.INIT_RAM_3E = 256'hFF3FFDFFFFFFFF9FFFFFFF7FFFFE0107FFFFFFFFFFFFFFF959FFFFFFFC7FFBFF;
defparam sdpb_inst_5.INIT_RAM_3F = 256'h997FFFFFFF9FFCFFFFFFFFDBFFFFFFC7FFFFC828FFFFFFFFFFFFFFFCB6FFFFFF;

SDPB sdpb_inst_6 (
    .DO({sdpb_inst_6_dout_w[30:0],sdpb_inst_6_dout[6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[6]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_6.READ_MODE = 1'b1;
defparam sdpb_inst_6.BIT_WIDTH_0 = 1;
defparam sdpb_inst_6.BIT_WIDTH_1 = 1;
defparam sdpb_inst_6.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_6.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_6.RESET_MODE = "SYNC";
defparam sdpb_inst_6.INIT_RAM_00 = 256'h0000000000000000000000017FFFFFFFF000000000012301A000000000000002;
defparam sdpb_inst_6.INIT_RAM_01 = 256'hEF888000000000000000000000000001FFFC7FFFE380000001040800A4000000;
defparam sdpb_inst_6.INIT_RAM_02 = 256'h16FFFFFBD423C880000000000000000000000001FFF9FFFFFF93112400B9FFA7;
defparam sdpb_inst_6.INIT_RAM_03 = 256'hFFFEC41BD3FFF7FFF7DADC00000000000000000000000000BFFDFFFFFFF2507A;
defparam sdpb_inst_6.INIT_RAM_04 = 256'hFFFE1FE37FFEFE4F7DEFFFFFFFFCFE00000000000000000000000000FFFEFFEF;
defparam sdpb_inst_6.INIT_RAM_05 = 256'h000000007F7EE1E3F7FDBA41D7CFFFFFFF878E06000000000000000000000000;
defparam sdpb_inst_6.INIT_RAM_06 = 256'h000000000000000001FC7E11FF7F8F200BBFFDEFFFFDDE500000000000000000;
defparam sdpb_inst_6.INIT_RAM_07 = 256'h08000000000000000000000001FF7FE1FFC00948013CFF7FFDFFFFE980000000;
defparam sdpb_inst_6.INIT_RAM_08 = 256'hF7BFFFE100000000000000000000000000EF3FF81FE38000009FFFAFAFFFEFF2;
defparam sdpb_inst_6.INIT_RAM_09 = 256'h0001FFFF3F7FFFFAC68000000000000000000000003783F8E1E3F8000003FFF7;
defparam sdpb_inst_6.INIT_RAM_0A = 256'h7FE0FFC00004FFF81CBFE7EFF020000000000000000000000017FC3C7E01FF00;
defparam sdpb_inst_6.INIT_RAM_0B = 256'h00009FFC3FF80FE600017DFC3C9FFFFFEC020000000000000000000000001FC0;
defparam sdpb_inst_6.INIT_RAM_0C = 256'h0000000000002FFE03F871E080003FFC7F73FFFFFF0100001020000000000000;
defparam sdpb_inst_6.INIT_RAM_0D = 256'h4000000000000000000000FE1CBC7F0020000BFF3F0E5FFFFF80E20900000000;
defparam sdpb_inst_6.INIT_RAM_0E = 256'hFFFE1C62018C0000000000000000018F1FC03FF1080006FF8E3413FFFFB50001;
defparam sdpb_inst_6.INIT_RAM_0F = 256'hF038008DFF7FF2090920000000000000000000080FFC3FFC020000FFE1B802FF;
defparam sdpb_inst_6.INIT_RAM_10 = 256'h00000007FE000021FF9BFFD440A0040000000000000000088FFF03FC0000003F;
defparam sdpb_inst_6.INIT_RAM_11 = 256'h011F8FC20010000CBF40037C3FFFEFED01408000000000000000000011FF183E;
defparam sdpb_inst_6.INIT_RAM_12 = 256'h0000000000818FFC206000009FD003E7CBFF7FE2A0010E000000000000000000;
defparam sdpb_inst_6.INIT_RAM_13 = 256'h3900000000000000002007FF800000000400006EF8FFFFEFC043293E4E000000;
defparam sdpb_inst_6.INIT_RAM_14 = 256'hAF090E2842E000000000000000D201FF980000000000002ED71FFFFE35944588;
defparam sdpb_inst_6.INIT_RAM_15 = 256'hFDE47FFFFD00005CC8000000000000000004001FC208000000008005E8E3FFFF;
defparam sdpb_inst_6.INIT_RAM_16 = 256'h000800081EEF87FFFFB4100140400000000000000000D081C000000000008100;
defparam sdpb_inst_6.INIT_RAM_17 = 256'h020485800000080083DCF0BFFFF8812026000000000000000001002004081000;
defparam sdpb_inst_6.INIT_RAM_18 = 256'h000004000081008000001C30007E9E0FFFFE00065BC400000000000000000240;
defparam sdpb_inst_6.INIT_RAM_19 = 256'h000000020080034010004080000008018007DEC0FFF900001BC0020000000000;
defparam sdpb_inst_6.INIT_RAM_1A = 256'h000C4A40000000000000000000009040800004000820FEF80AF78800C5EACA00;
defparam sdpb_inst_6.INIT_RAM_1B = 256'h778AAC00002EEC200000000000000000410000384000220000841FCF80BFF800;
defparam sdpb_inst_6.INIT_RAM_1C = 256'h0002007CF0006028019E54A000000008220404000083510220000800000003ED;
defparam sdpb_inst_6.INIT_RAM_1D = 256'h000000100000000FF020100006A9AA8400000000200000008800001000000000;
defparam sdpb_inst_6.INIT_RAM_1E = 256'h002201030800002000001001F04000000239ABA1800000008045040000201008;
defparam sdpb_inst_6.INIT_RAM_1F = 256'h0000000000184004440000000000040020000000000020364000000004000040;
defparam sdpb_inst_6.INIT_RAM_20 = 256'h7000000000080000000104020000000200000000040000000100793640000000;
defparam sdpb_inst_6.INIT_RAM_21 = 256'h2008091845000000000000008000101888000000400000000100000000001F83;
defparam sdpb_inst_6.INIT_RAM_22 = 256'h0010000000003B6B4EE000000000000000000180410000001080004000600000;
defparam sdpb_inst_6.INIT_RAM_23 = 256'h000000008006000000001031BD80000000000000000000004080000002000001;
defparam sdpb_inst_6.INIT_RAM_24 = 256'h000000000010800040018000000002401A860000000000000080000010000000;
defparam sdpb_inst_6.INIT_RAM_25 = 256'h00040000026000000002050060002000000000034B0100000000000000000000;
defparam sdpb_inst_6.INIT_RAM_26 = 256'h0000000000000000000000000000800040000C00000000060A46600000000000;
defparam sdpb_inst_6.INIT_RAM_27 = 256'h223FC00000000000400080000000000000000C02400001800002000A08444000;
defparam sdpb_inst_6.INIT_RAM_28 = 256'h00000000072FD8000000000000003000000000000000009BC000003000000008;
defparam sdpb_inst_6.INIT_RAM_29 = 256'h00000000C000780003CEFE000000000002005C00000000000000000000000006;
defparam sdpb_inst_6.INIT_RAM_2A = 256'h0000000000004C001E007F00000D4F38000000000011FF000000000000000000;
defparam sdpb_inst_6.INIT_RAM_2B = 256'h00000000000000000000000000F27FE0010C3C70000000000003FF8000000000;
defparam sdpb_inst_6.INIT_RAM_2C = 256'h000005E000000000000000000000008000013F7C0109880700000000000028E0;
defparam sdpb_inst_6.INIT_RAM_2D = 256'h00000000000000C000000000000000000000004000003F7B805E0A1F00000000;
defparam sdpb_inst_6.INIT_RAM_2E = 256'hAE020061A900000000000000000000000000000000000100000005F9D0001047;
defparam sdpb_inst_6.INIT_RAM_2F = 256'h0000001FADC000192000000000000000000000000000000000000000000000B7;
defparam sdpb_inst_6.INIT_RAM_30 = 256'h0000780000000003FCF810025200000000000000004000000000000000000FC0;
defparam sdpb_inst_6.INIT_RAM_31 = 256'h04200000000FC000000000007EF704090D400000000000000018800000000000;
defparam sdpb_inst_6.INIT_RAM_32 = 256'h000200000000800003E00000000000000FF3E08004A000000000000000058000;
defparam sdpb_inst_6.INIT_RAM_33 = 256'h0000000000018A00000000000F0000000000000001EFDC20000A000000000000;
defparam sdpb_inst_6.INIT_RAM_34 = 256'h882100000000000000004580000002001C00000000001C00003F5B0002084000;
defparam sdpb_inst_6.INIT_RAM_35 = 256'h0000F9EC0080180000000000000048C00000008038000000000001000007F9E0;
defparam sdpb_inst_6.INIT_RAM_36 = 256'h0000000000001FE7800138000000000000000860000000003000000600000800;
defparam sdpb_inst_6.INIT_RAM_37 = 256'h2000028000000000000003EF3000180000000000000000300001000020000040;
defparam sdpb_inst_6.INIT_RAM_38 = 256'h0000080020000000000000000024007EBA000000000000000000001000000000;
defparam sdpb_inst_6.INIT_RAM_39 = 256'h000000060000000430000500000000000004000EB5C018800000000000000208;
defparam sdpb_inst_6.INIT_RAM_3A = 256'h000000000000000100000004100000000000000000000001F2DC002100000000;
defparam sdpb_inst_6.INIT_RAM_3B = 256'h07CA70020000000000000000800000001800020000000000000010003BCF8010;
defparam sdpb_inst_6.INIT_RAM_3C = 256'h0000000000FF3A008C000000000000006000000008000A000000000000000000;
defparam sdpb_inst_6.INIT_RAM_3D = 256'h0000000000000000001F79C00000000000000008300000000600020000000000;
defparam sdpb_inst_6.INIT_RAM_3E = 256'h0080000000000000000000000003FCF800000000000000000800000001000200;
defparam sdpb_inst_6.INIT_RAM_3F = 256'h03000000004000000000000000000000000075D7000000000000000006000000;

SDPB sdpb_inst_7 (
    .DO({sdpb_inst_7_dout_w[30:0],sdpb_inst_7_dout[7]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_7.READ_MODE = 1'b1;
defparam sdpb_inst_7.BIT_WIDTH_0 = 1;
defparam sdpb_inst_7.BIT_WIDTH_1 = 1;
defparam sdpb_inst_7.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_7.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_7.RESET_MODE = "SYNC";
defparam sdpb_inst_7.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC;
defparam sdpb_inst_7.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00FFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_04 = 256'hFFFFE01CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF001F;
defparam sdpb_inst_7.INIT_RAM_05 = 256'hFFFFFFFFFFFF1E1C0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFF81EE00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF801E003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC007E01C7FFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC071E1C07FFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0A = 256'h801F003FFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC3C381FE00FF;
defparam sdpb_inst_7.INIT_RAM_0B = 256'hFFFFE003C007F019FFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE03F;
defparam sdpb_inst_7.INIT_RAM_0C = 256'hFFFFFFFFFFFFF001FC078E1C7FFFFFFF808FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFF01E3C380FE1FFFFFFFC0F1FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE70E03FC00E07FFFFFFF1C00FFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_0F = 256'hFFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7F003C00381FFFFFFFE4001FF;
defparam sdpb_inst_7.INIT_RAM_10 = 256'h887FFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07000FC03A0FFFFFF;
defparam sdpb_inst_7.INIT_RAM_11 = 256'h82E0703DC227FFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0E00E7C1;
defparam sdpb_inst_7.INIT_RAM_12 = 256'hFFFFFFFFF04E7003C091FFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFF10F80070387FFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF240E00640C1FFFFFFFFFC000FFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_15 = 256'h0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE383E0310607FFFFFF7FF8001FFFFF;
defparam sdpb_inst_7.INIT_RAM_16 = 256'hFFF00007E0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8204E384683FFFFF808FF;
defparam sdpb_inst_7.INIT_RAM_17 = 256'h0C03081FFFFC00017C000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0E10F813217F;
defparam sdpb_inst_7.INIT_RAM_18 = 256'hFFFFF84781008307FFFC03C00F8001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC126;
defparam sdpb_inst_7.INIT_RAM_19 = 256'hFFFFFFF9F0FFFC986060A041FFFF07FE01F8003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFC3C3C7F9E0E1848307FFF83FFF01F0007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1B = 256'h087FFFFFFFFFFFFFFFFFFFFF0F0F0FE182E666043FFFC1FFFF03E0007FFFFFFF;
defparam sdpb_inst_7.INIT_RAM_1C = 256'hFFFC1F800001FFFFFFFFFFFFFFFFFFF0C1F3C3FC384CA0911FFFF0FFFFE07C00;
defparam sdpb_inst_7.INIT_RAM_1D = 256'h1FFFFF0FFFFF87F000000FFFFFFFFFFFFFFFFFFC1E3CF3FF0590F0285FFFFC3F;
defparam sdpb_inst_7.INIT_RAM_1E = 256'hFF41820407FFFFC3FFFFE0FE000001FFFFFFFFFFFFFFFFFF038200FFF11C0804;
defparam sdpb_inst_7.INIT_RAM_1F = 256'hFF80001FFFE030C283FFFFF0FFFFF87FC000003FFFFFFFFFFFFFFFFFF800003F;
defparam sdpb_inst_7.INIT_RAM_20 = 256'hFFFFFFFFFFF00007FFFE0B3133FFFFFC1FFFFE1FF8000007FFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_21 = 256'h1FFFFFFFFFFFFFFFFFFF00007FFFE32505FFFFFF83FFFF07FE000000FFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_22 = 256'hFFE0000007FFFFFFFFFFFFFFFFFFFC001FFFFE4380FFFFFFE07FFF83FF800000;
defparam sdpb_inst_7.INIT_RAM_23 = 256'hFF87FFC07FF8000001FFFFFFFFFFFFFFFFFFFE0003FFFFF0207FFFFFFC1FFFC0;
defparam sdpb_inst_7.INIT_RAM_24 = 256'hE23FFFFFFFE07FE03FFE0000007FFFFFFFFFFFFFFFFFFF80007FFFFE087FFFFF;
defparam sdpb_inst_7.INIT_RAM_25 = 256'h0003FFFFFC9FFFFFFFFC02401FFFC000001FFFFFFFFFFFFFFFFFFFE0001FFFFF;
defparam sdpb_inst_7.INIT_RAM_26 = 256'hFFFFFFFE0001FFFFFFFFFFFFFFFF00003FFFF0000007FFFFFFFFFFFFFFFFFFF8;
defparam sdpb_inst_7.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFF80007FFFFFFFFFFFFFFFF0003FFFFE000001FFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_28 = 256'h00003FFFFFFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFFFFF003FFFFFC00000FFFF;
defparam sdpb_inst_7.INIT_RAM_29 = 256'hFFFFFFFF000007FFFFFFFFFFFFFFFFFFFC0003FFFFFFFFFFFFFFFFFFFFFFFFF8;
defparam sdpb_inst_7.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFE00000FFFFFFFFFFFFFFFFFFFFE000FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF00001FFFFFFFFFFFFFFFFFFFFC007FFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2C = 256'hFFFFF81FFFFFFFFFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFFFC01F;
defparam sdpb_inst_7.INIT_RAM_2D = 256'hFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2E = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE3FFFFFF8000FFFFFFF;
defparam sdpb_inst_7.INIT_RAM_2F = 256'hFFFFFFE0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0FFFFFFF00;
defparam sdpb_inst_7.INIT_RAM_30 = 256'hFFFF87FFFFFFFFFC0007FFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFFFFFFFFF03F;
defparam sdpb_inst_7.INIT_RAM_31 = 256'hF81FFFFFFFF03FFFFFFFFFFF8000FFFFFFFFFFFFFFFFFFFFFFC07FFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_32 = 256'hFFF847FFFC007FFFFC1FFFFFFFFFFFFFF0001FFFFFFFFFFFFFFFFFFFFFE01FFF;
defparam sdpb_inst_7.INIT_RAM_33 = 256'hFFFFFFFFFFFC21FFFE000FFFF0FFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFF107FFF8001FFE3FFFFFFFFFFE3FFFFC000FFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_35 = 256'hFFFF0003FFFFFFFFFFFFFFFFFFFF803FFFE0007FC7FFFFFC000000FFFFF8001F;
defparam sdpb_inst_7.INIT_RAM_36 = 256'hFFFFFFFFFFFFE0007FFFFFFFFFFFFFFFFFFFE01FFFF8003FCFFFFF81FFFFF7FF;
defparam sdpb_inst_7.INIT_RAM_37 = 256'hDFFFFC7FFFFFFFFFFFFFFC000FFFFFFFFFFFFFFFFFFFF00FFFFE001FDFFFFE3F;
defparam sdpb_inst_7.INIT_RAM_38 = 256'hFFFFF007DFFFFCFFFFFFFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFF80FFFFFC00F;
defparam sdpb_inst_7.INIT_RAM_39 = 256'hFFFFFF01FFFFFE03CFFFF8FFFFFFFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFC07;
defparam sdpb_inst_7.INIT_RAM_3A = 256'hFFFFFFFFFFFFFF80FFFFFFC3EFFFF9FFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3B = 256'hF8000FFFFFFFFFFFFFFFFFC07FFFFFFFE7FFF9FFFFFFFFFFFFFFFFFFC0007FFF;
defparam sdpb_inst_7.INIT_RAM_3C = 256'hFFFFFFFFFF0001FFFFFFFFFFFFFFFFE01FFFFFFFF7FFF1FFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFF00FFFFFFFF9FFF9FFFFFFFFFF;
defparam sdpb_inst_7.INIT_RAM_3E = 256'hFF7FFDFFFFFFFFFFFFFFFFFFFFFC0007FFFFFFFFFFFFFFFC07FFFFFFFEFFF9FF;
defparam sdpb_inst_7.INIT_RAM_3F = 256'h00FFFFFFFFBFFEFFFFFFFFFFFFFFFFFFFFFF8000FFFFFFFFFFFFFFFE01FFFFFF;

SDPB sdpb_inst_8 (
    .DO({sdpb_inst_8_dout_w[29:0],sdpb_inst_8_dout[1:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_8.READ_MODE = 1'b1;
defparam sdpb_inst_8.BIT_WIDTH_0 = 2;
defparam sdpb_inst_8.BIT_WIDTH_1 = 2;
defparam sdpb_inst_8.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_8.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_8.RESET_MODE = "SYNC";
defparam sdpb_inst_8.INIT_RAM_00 = 256'h9FEFF0DFD5140FF84104040EB6EDB2F01905BE954C6A400FDCEBF3BFFE29D370;
defparam sdpb_inst_8.INIT_RAM_01 = 256'hFFCB3FBCCCFBA4883948743B2985AAADA654436418FF816A6BAB8FFFC0002121;
defparam sdpb_inst_8.INIT_RAM_02 = 256'h5595ABFFFB1C0356DEBECFFEC34403D5FF3555413FF761EF6F8C065961DAB30B;
defparam sdpb_inst_8.INIT_RAM_03 = 256'hAD31FC55B4CC66EF6F0BAFAA0BEDA93EC9204829B15565AC4AA82B35C17A90C5;
defparam sdpb_inst_8.INIT_RAM_04 = 256'h56A5F8FA2033A3C01046A9AABF801CB9F3E7EFEF31B3200A39BC3443C332E15E;
defparam sdpb_inst_8.INIT_RAM_05 = 256'h78892FF030B8BC05D15757A01460F9868FF29EEAAEFB9D77ACAD85CCE8466156;
defparam sdpb_inst_8.INIT_RAM_06 = 256'hA5C9421292CD555159114F51B43E4A46DD29496ABEAFBC3350EA3ABFEFFC3F0F;
defparam sdpb_inst_8.INIT_RAM_07 = 256'hF5CCC0BF3CFFF8CF3285DBF0F0B31F64D973649D8C452F5AAFFC8ABEAEA8A62C;
defparam sdpb_inst_8.INIT_RAM_08 = 256'h1FBAFFE68DB5955F0DA36B10776C4546554414ED69BFE8A4F2D95596AAABAF03;
defparam sdpb_inst_8.INIT_RAM_09 = 256'h2715515465ABBAF330EA792CF3FFCFF3FCF2369FC3FFEABB9C2153E4EAC00002;
defparam sdpb_inst_8.INIT_RAM_0A = 256'hA50768C1828BC0C917BCCF3EEF6A956C8D39F754B946015159551009282FF85B;
defparam sdpb_inst_8.INIT_RAM_0B = 256'h155551CEFF7AFA04EB7010F111A59AAAEF0F0D121BFFF3BF3FFF5628AFF3FAAA;
defparam sdpb_inst_8.INIT_RAM_0C = 256'hFFFFFFBC2FFFE86AA98389085F977BC2C4A2CFC2EAB955CDB091AA10F3E4A305;
defparam sdpb_inst_8.INIT_RAM_0D = 256'hB6C3F490638246F341FD44428FE9FF8A56DB3365F0455566AFF8CEC65D7FFF0F;
defparam sdpb_inst_8.INIT_RAM_0E = 256'h69B6C0FBCF16F030CF3C39D8623FFDEAB5590E9642601C63BD0AAFCEF9A65D64;
defparam sdpb_inst_8.INIT_RAM_0F = 256'hEFD08EFFEBFAA4FA2ED27DABCBF7A718041C140031031FE7E6C2B0C0C00D5655;
defparam sdpb_inst_8.INIT_RAM_10 = 256'hC89628FFF33040505556AEBF23489FB0FF3F2AAA7566BBABAA6644229E2FB44A;
defparam sdpb_inst_8.INIT_RAM_11 = 256'h659940008D2072EC69941B7FFEEA6D796F1CEF58C26B9CB1B010FC000ED176A9;
defparam sdpb_inst_8.INIT_RAM_12 = 256'hCABF0003C396B3A6458C22AFFF03F3001055D5AA8F6EF38167DB56427666AAA6;
defparam sdpb_inst_8.INIT_RAM_13 = 256'h0C0CDFB4359795A2A89254413E59BB137AE575AAABAEBA721104780AD233AFAA;
defparam sdpb_inst_8.INIT_RAM_14 = 256'h4C9412F6AF0CCF38296FFFCFFFA866D956F03B5EFEC03FFF333FB14065935BCC;
defparam sdpb_inst_8.INIT_RAM_15 = 256'hFFFBFABEFDFEEE52B31F12A3EA88D6569505457CF0F490583506CF4D9AE3A99B;
defparam sdpb_inst_8.INIT_RAM_16 = 256'h28267F7C6AABAAA5BB5C68A311B51F9451CAFCF0EFC920D5938028D5BFCFFFFF;
defparam sdpb_inst_8.INIT_RAM_17 = 256'h5532A3AB5FBFCFFAAFFA65A2551F32573C676276B2C23159276404504FCFCB72;
defparam sdpb_inst_8.INIT_RAM_18 = 256'h9045101040B8FF857DCCF9CB017BBBE8120087A907C4E64E174C57FAFEEBDDA4;
defparam sdpb_inst_8.INIT_RAM_19 = 256'hA030C66BFB3BA44285590869B1ABAFBBCA869570398D11560C3165AA69CCB805;
defparam sdpb_inst_8.INIT_RAM_1A = 256'hE6D436F81511A6B011D404000CBEDEF935155D587256A6A720BEE71A920FF8F5;
defparam sdpb_inst_8.INIT_RAM_1B = 256'h40E74460818B0B04100CA867AFAEA984E8079AC798125AAEBA58040F13A595BA;
defparam sdpb_inst_8.INIT_RAM_1C = 256'h69654C3D7E4742C8C1B4AFC2D3F15157B154F3FCA273AFEA9BD43222C305AAA9;
defparam sdpb_inst_8.INIT_RAM_1D = 256'hAE5C455683FF55661541823B15A074DE80A0436DABDEE95BA4CFE470EDBF5525;
defparam sdpb_inst_8.INIT_RAM_1E = 256'h67903E335EEB3597D08A5FCED34E6BF2C5038DF2C0BF01429EC03FDEBEEBBAAF;
defparam sdpb_inst_8.INIT_RAM_1F = 256'h15AB0EEFAFEEA9FADAFD08AA83C00496514E1DBDB8668DC84E0B269B5A69B99D;
defparam sdpb_inst_8.INIT_RAM_20 = 256'hCF4A26FDF05555950BB1FE92DCD2AC1555590438949DBBADE3BDADEF9F15AFC4;
defparam sdpb_inst_8.INIT_RAM_21 = 256'h94A95EBCDC1B256F055BB3BBA9BE9BA6AE6BE90FAC7CE045554FEF7419C4CC3A;
defparam sdpb_inst_8.INIT_RAM_22 = 256'h044F88672B7C81D242D41589CB15595910DC2EA517521BCC1641D503A426E54D;
defparam sdpb_inst_8.INIT_RAM_23 = 256'h114110031939C51895CC737BCC0A1C55BCD556FBEAAE6ABAEA6EF66B167B1687;
defparam sdpb_inst_8.INIT_RAM_24 = 256'hA651AA9AA70EA91AFF0F9DBAB9C46747D3BB01343080D641940A1BF9C8732243;
defparam sdpb_inst_8.INIT_RAM_25 = 256'h200042EB5C833E04F0C0000F0F4E71C4E6013FDE95FD5D4D6AB0056ACA99AA5A;
defparam sdpb_inst_8.INIT_RAM_26 = 256'h4559F045A2AA9A9558999566A9653D35A8CB998A800DA8481A277581E7587459;
defparam sdpb_inst_8.INIT_RAM_27 = 256'h4ACE68BFDD850D004F0CE24A9508C1115B00C03F3E5748560A3B6221FD24ACB7;
defparam sdpb_inst_8.INIT_RAM_28 = 256'hB5AD1DD35730B55A2D56A6B1042965695154055555614253D9BAA687E07350E4;
defparam sdpb_inst_8.INIT_RAM_29 = 256'h315A97F011FAE655EB4E7B74261C6A3C003C3A13994FA01ED5ACF33EFAA43759;
defparam sdpb_inst_8.INIT_RAM_2A = 256'hDD66ABCFFEF93DDB9581DD822378743DCCD1C95AF005A654E401544016196013;
defparam sdpb_inst_8.INIT_RAM_2B = 256'h54CC430340031D200ED198EE0590FA1C942CF011E5E32498107003A6C417E1D9;
defparam sdpb_inst_8.INIT_RAM_2C = 256'hBAE0BCA1162F6F37DE15A6FBAEA4FE9B0B565ABE31E8F4AE1179C6992BFFC551;
defparam sdpb_inst_8.INIT_RAM_2D = 256'hF5F00AFE8E459FC307F3100F0C044F0307FD453AD6B86FFC0440C703A124756F;
defparam sdpb_inst_8.INIT_RAM_2E = 256'h89AA1C06468B44D17BB6FFA99471474A34EC1EB79AAA42922B9E9AFEB1170E33;
defparam sdpb_inst_8.INIT_RAM_2F = 256'h9DA22739541D624380D7BF6FDB15417C34FF1CBA30F32322F36DF71F84FE65D8;
defparam sdpb_inst_8.INIT_RAM_30 = 256'h3F24A8BEB4A70AC72D10F001C5C01BF189EEAEAD0B7F6B9F3D63FC6A7B39533A;
defparam sdpb_inst_8.INIT_RAM_31 = 256'h2BCE1FD26A5541F86FB8160B59BB8A500462D65A01D201466F8F6F2BEFBDEBBE;
defparam sdpb_inst_8.INIT_RAM_32 = 256'h45655956BCEAAAAFE7A8DE5C371BAAA3639A10F4266A898C0B5E96BB83221C29;
defparam sdpb_inst_8.INIT_RAM_33 = 256'hC05559A5A7E0F4B2CC328DBC5E64244F93B6D644B4A573687928DAE81075B201;
defparam sdpb_inst_8.INIT_RAM_34 = 256'h293FC409C58569C6F4FF5550156A9997E69AAA473929CAD12BCEC020450686A9;
defparam sdpb_inst_8.INIT_RAM_35 = 256'h546569E550AC1C421FC004185504DCE74071FF0A0042D14EEB071A887E6B69B8;
defparam sdpb_inst_8.INIT_RAM_36 = 256'h3A5E33B7E4BFBE12FCFFE5815F20018346A900555402AE9A9C95915D4391CD71;
defparam sdpb_inst_8.INIT_RAM_37 = 256'hA5065511F229D8A735A569AAA92A501312F70100173DB8E5BFA2C471AC051040;
defparam sdpb_inst_8.INIT_RAM_38 = 256'h77B9EA57CAC013003B94231C960AD0361162720E1AE05D30DE0B2BFB35107564;
defparam sdpb_inst_8.INIT_RAM_39 = 256'hD576282A73005CC15456500D6807B19FF4ABFDF6BE369E06BA5BF083CCF8D767;
defparam sdpb_inst_8.INIT_RAM_3A = 256'h0EF5BFC933DCB931DF9A4F097168B00CCBEACE76592A33206D38CB6AAD08BACC;
defparam sdpb_inst_8.INIT_RAM_3B = 256'h11BE2AD238D12A04676C898BA9BF000F00D4313C5ADBF55EEAC6C33FFFCBCDB0;
defparam sdpb_inst_8.INIT_RAM_3C = 256'h027783940F30189BE0240BEFEFFEA64DE8B59342BA0AAE33CBAE6038BFAF887E;
defparam sdpb_inst_8.INIT_RAM_3D = 256'hEFFAA64E97164FD986591E11AE6388FDC6772CB7B956E3000F03000C8C2CBE0E;
defparam sdpb_inst_8.INIT_RAM_3E = 256'h7F830273FFF2F2AC258D7E0566D32FF6807B86BFB9BFEA9397BC07929DA155DB;
defparam sdpb_inst_8.INIT_RAM_3F = 256'hF63EAC25F45916AAA2BFA540E5DEAD543B2C1E0BDE78E189CA0FBAC849ED45EE;

SDPB sdpb_inst_9 (
    .DO({sdpb_inst_9_dout_w[29:0],sdpb_inst_9_dout[3:2]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_9.READ_MODE = 1'b1;
defparam sdpb_inst_9.BIT_WIDTH_0 = 2;
defparam sdpb_inst_9.BIT_WIDTH_1 = 2;
defparam sdpb_inst_9.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_9.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_9.RESET_MODE = "SYNC";
defparam sdpb_inst_9.INIT_RAM_00 = 256'h6AAAAFBABFFFF9AC2FFFFFFAA8855EC56AFFFFFFF955AAA5665559555595543E;
defparam sdpb_inst_9.INIT_RAM_01 = 256'h556595566655550F9A042EF05555555555553571550CB155555565556AAA96F1;
defparam sdpb_inst_9.INIT_RAM_02 = 256'h5555555555A6A9421EAABAAABEFFFEA763EFFFFFEAA11C16D567FFFFFF9559A5;
defparam sdpb_inst_9.INIT_RAM_03 = 256'h15B55BFFFFB9555595A555559555554FA351A26C0555555555554DBC1543D715;
defparam sdpb_inst_9.INIT_RAM_04 = 256'h555500CB0544DA8555555555556AA655B2CAAAAAEEAEEFFABB5FEFFEBEEE4855;
defparam sdpb_inst_9.INIT_RAM_05 = 256'hE9FC2AAFEFABAA41D5415D6FFFFF85656559555555555543E78D1E07C1555555;
defparam sdpb_inst_9.INIT_RAM_06 = 256'hE99CD87DB01155555555501CB14005DC1155555555555699502CAAAAAAABEAFA;
defparam sdpb_inst_9.INIT_RAM_07 = 256'h5528CAAAEBAAABBAEEAF2AAFAFAEEAA9C5511554BBFFE8555556655555565550;
defparam sdpb_inst_9.INIT_RAM_08 = 256'h5555555565555553E51D85665B015555555555359C000E2FC5155555555555A9;
defparam sdpb_inst_9.INIT_RAM_09 = 256'hB0555555555555599A576F2BAEAABAAEABA926DABEAAAAAAA3115495D6BFFFD5;
defparam sdpb_inst_9.INIT_RAM_0A = 256'hAA9755D505BABFB955566595555555409022AA5F36C0555555555553AF000088;
defparam sdpb_inst_9.INIT_RAM_0B = 256'h55555510D8B000368F0555055555555555A55B8BAAAAAEAAEAAA9C5AAAAEAAAA;
defparam sdpb_inst_9.INIT_RAM_0C = 256'hAAAAA4322AAAABAAAAA90D517459DABE915965695555550FC0EE1B652C6C0455;
defparam sdpb_inst_9.INIT_RAM_0D = 256'h30C3AE7560DAC00455015554081C000E2EC044450555555555566536BEAAAAFA;
defparam sdpb_inst_9.INIT_RAM_0E = 256'h55556A54A902AFEFBAEBEA615AEAAAAAAAAAA435E51456AEA955556555555140;
defparam sdpb_inst_9.INIT_RAM_0F = 256'hAA955555555555033C00DB862C5C6F015551555543BE0003A140051515515555;
defparam sdpb_inst_9.INIT_RAM_10 = 256'hF60B0100044555555555555597A6FAAFAAEAEA4C1BAAAAAAAAAAAA91D0514662;
defparam sdpb_inst_9.INIT_RAM_11 = 256'hAAAAAAAA434185317AA9555555555540FC0CFB4C30D882B00555015550E6B000;
defparam sdpb_inst_9.INIT_RAM_12 = 256'hC0005554140CFF000E8AF0000054045555551555654B9CD6AAAAA95C145AAAAA;
defparam sdpb_inst_9.INIT_RAM_13 = 256'hFA6A64EF7325AAAAAAAAAAAA95DD00501D9A8555555555443500EE3F8304221B;
defparam sdpb_inst_9.INIT_RAM_14 = 256'h0E803C036ED01D4DBC00001000009AC003896F00001540004440055555543117;
defparam sdpb_inst_9.INIT_RAM_15 = 256'h00000000010000D837BAFFECEA096AAAAAAAAA965A5775694403645555595554;
defparam sdpb_inst_9.INIT_RAM_16 = 256'h300049815555555503A00FDAF09C50138BC00105001038F003F837C000100000;
defparam sdpb_inst_9.INIT_RAM_17 = 256'h003E54BF0000100000000000000F1003CBA3CE6E5B505AAAA9AAAAAAA5655DC4;
defparam sdpb_inst_9.INIT_RAM_18 = 256'hAAAAAAAAAA56557747903024555555555439C38FFFF8F012777C000000000EF8;
defparam sdpb_inst_9.INIT_RAM_19 = 256'h113BC000004000DEC00FECDBF0000000100000303FFAC0AB8CE891119D3156AA;
defparam sdpb_inst_9.INIT_RAM_1A = 256'hA99C3F969B05555AAA6AAAAAA6556555DD036C0185555554553E1FF67FFBDC01;
defparam sdpb_inst_9.INIT_RAM_1B = 256'h5503E8EF57FF4C01911CAC000000000EDC03F951BC0000000000000F3EA904EA;
defparam sdpb_inst_9.INIT_RAM_1C = 256'h00000C3FEAA439AFBEAADBC3C00555555AAA5956595955555225684410555555;
defparam sdpb_inst_9.INIT_RAM_1D = 256'h55599000158055555554F289F13260B06A575AFC000000039BCFFF8E2BFF0000;
defparam sdpb_inst_9.INIT_RAM_1E = 256'h35F03FE8B6BF3000C0000FCFFEA53A2B4FF8A0DFC0005555556A956555555555;
defparam sdpb_inst_9.INIT_RAM_1F = 256'h5555A555555555555555BB401421555555500334EFF8AEE556D1ADBF0000000C;
defparam sdpb_inst_9.INIT_RAM_20 = 256'h11CDB11BF000000003FBFFFE746FFC000000003FFFA538EAB92E6A4C3F000015;
defparam sdpb_inst_9.INIT_RAM_21 = 256'h86542FAA3F7F000055555955555555555555551C41570555555000BD7CC3564B;
defparam sdpb_inst_9.INIT_RAM_22 = 256'h55501B7DCF2C03C3157B9706BF00000000F7BFFFE7CAFFCC0000C003FFE90E19;
defparam sdpb_inst_9.INIT_RAM_23 = 256'h000000033FEA538684A68872B9293C00011555555555555555555554F1D48414;
defparam sdpb_inst_9.INIT_RAM_24 = 256'h55555555543BC14000500F8AE0BC0067C4585EFDAFC0C000000EABFFFA5CAFC3;
defparam sdpb_inst_9.INIT_RAM_25 = 256'h0000D6BFFBA5C6FCF0C0000F0FFA94A1E9AA97A157E74ACC0005555565555555;
defparam sdpb_inst_9.INIT_RAM_26 = 256'hC000055559555555555555555555414401100EA7F0073060005582E31AFC3000;
defparam sdpb_inst_9.INIT_RAM_27 = 256'h8FD1754786BF0C000F0CFE8BFFFA2DAFFF00C03F3FFEA538A6C6A99A4214A2EE;
defparam sdpb_inst_9.INIT_RAM_28 = 256'h26A1FB79A99FC0956E000005555555555555555555555554000003254DF73CC3;
defparam sdpb_inst_9.INIT_RAM_29 = 256'h440003C694FF35ECE0FB028DA1ABFF3C003C3F97BFFA9ED6BFFCF33FFFFFE94E;
defparam sdpb_inst_9.INIT_RAM_2A = 256'h6BFFFFCFFFFFEA539F1EABABAB5691878149C000055555551555555555555554;
defparam sdpb_inst_9.INIT_RAM_2B = 256'h5511545455545145500000F75531FFDE87CE842F731AFFFC003003E4CBFEA98D;
defparam sdpb_inst_9.INIT_RAM_2C = 256'hFFF0FCFE08AAE989D6FFFFFFFFFFAAA43763AFEEEA4646537FE36AC000001555;
defparam sdpb_inst_9.INIT_RAM_2D = 256'h115B961BC000001454045550515550545400003E0C2C4CFCBC70C336ED76AFFF;
defparam sdpb_inst_9.INIT_RAM_2E = 256'hC0200C0BECD76BBFFFFFFFFFA50ABAA4916BFFFFFFFFFEA94D2D81FFDAA9A398;
defparam sdpb_inst_9.INIT_RAM_2F = 256'h50DF81EA3EA6AAA9BA6B9B9C8B00000145005100450444440440330F9F834480;
defparam sdpb_inst_9.INIT_RAM_30 = 256'h404100FFE82F1160000DF0007EA285AFFFFFFFFFF9E06AA5461AABFFFFFFFEEA;
defparam sdpb_inst_9.INIT_RAM_31 = 256'h91F1AABFFFFFFFAA9439992EFA955A8AAA96AAAFB6FB00000010000000000000;
defparam sdpb_inst_9.INIT_RAM_32 = 256'h00000000010000000001000C3EAAFF80000198F00588286BFFFFFFFFFE9886AA;
defparam sdpb_inst_9.INIT_RAM_33 = 256'hBFFFFFFFFEA9995A651326ABFFFFFFFAA9434187F0CF32A8A9A9BEEBA0B0EF00;
defparam sdpb_inst_9.INIT_RAM_34 = 256'hAABA600FFFA1202FFCFF000000000003000000033FE57FC0401156600064B686;
defparam sdpb_inst_9.INIT_RAM_35 = 256'h0000001C0001E6BDAABFFFFFFFFA5C85AA4D31AAFFFFBFFAA9A437CA1F0E33CA;
defparam sdpb_inst_9.INIT_RAM_36 = 256'hEAA5426ED8FEF103CE56A4020F3FE1217BFF0000000000000000000C03FE6BF0;
defparam sdpb_inst_9.INIT_RAM_37 = 256'h00000000F33FA7FF300000000000548C1AAEFFFFFEEA940C5554F85AABFFFFFF;
defparam sdpb_inst_9.INIT_RAM_38 = 256'hC55536C56ABFFEFFEAAA9437F793BEE85C01A810C000FF953E2AFFFF30003000;
defparam sdpb_inst_9.INIT_RAM_39 = 256'h515CEAFFF3000CC00000000C3C0FEE4FB0000000000015C721AAAFBEBBABA97C;
defparam sdpb_inst_9.INIT_RAM_3A = 256'hAF1AAABBEEBBAA941C55528D5AABAFFBBAAA65438079A45AA8690DB5555100CA;
defparam sdpb_inst_9.INIT_RAM_3B = 256'h9AABF12C98595050E8BC7202FFFF000F00C0303C0FFFFFA45AC014400010143E;
defparam sdpb_inst_9.INIT_RAM_3C = 256'h901B1455504557B00E86AAAAAAAAAAA526C55425C5AAAAEEBAAAAA9538AB6769;
defparam sdpb_inst_9.INIT_RAM_3D = 256'hAAAAAAA553E1684148C2AA24301AA6500DA59C2BAFFFF3000F03000CCC3CFFFA;
defparam sdpb_inst_9.INIT_RAM_3E = 256'hFFC30333FFF3F3FFE9349881951455DB38CC6AAAAAAAAAA9511D540DAD5AAAAA;
defparam sdpb_inst_9.INIT_RAM_3F = 256'h54DDC1403315AAAAAEAAAAAA550E716EE7C5BA8E3F665A9550D77E9C346BFFFF;

SDPB sdpb_inst_10 (
    .DO({sdpb_inst_10_dout_w[29:0],sdpb_inst_10_dout[5:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_10.READ_MODE = 1'b1;
defparam sdpb_inst_10.BIT_WIDTH_0 = 2;
defparam sdpb_inst_10.BIT_WIDTH_1 = 2;
defparam sdpb_inst_10.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_10.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_10.RESET_MODE = "SYNC";
defparam sdpb_inst_10.INIT_RAM_00 = 256'hFFFFFFFFFFFFFF96BFFFFFFFFF80080303FFFFFFFFFFFFFFFFFFFFFFFFFFFFEA;
defparam sdpb_inst_10.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFA9584C6AFFFFFFFFFFFFFE0AFFFF95FFFFFFFFFFFFFFFFE5A;
defparam sdpb_inst_10.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFF9A7FFFFFFFFFFFFFD59FFFFFFFFFE0402800FFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_03 = 256'h84103FFFFFFFFFFFFFFFFFFFFFFFFFFAA9AA61ABFFFFFFFFFFFFF81BFFFE56FF;
defparam sdpb_inst_10.INIT_RAM_04 = 256'hFFFFFF26FFFFA4BFFFFFFFFFFFFFFFFF997FFFFFFFFFFFFFE5A7FFFFFFFFF803;
defparam sdpb_inst_10.INIT_RAM_05 = 256'hFF56FFFFFFFFFFF0801808FFFFFFFFFFFFFFFFFFFFFFFFFEA956D76ABFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_06 = 256'hAA2685C6AFFFFFFFFFFFFFE1AFFFF9EBFFFFFFFFFFFFFFFFFE56FFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_07 = 256'hFFE66FFFFFFFFFFFFFF9ABFFFFFFFFFF8028C103FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFEAA9D61A1AAFFFFFFFFFFFFE82BFFFAA6BFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_09 = 256'hAFFFFFFFFFFFFFFFFFFE55BFFFFFFFFFFFFFDABFFFFFFFFFFE0001404FFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0A = 256'hFFFF0240102FFFFFFFFFFFFFFFFFFFFFAA9757D75ABFFFFFFFFFFFFEB6FFFFA5;
defparam sdpb_inst_10.INIT_RAM_0B = 256'hFFFFFFFFA1AFFFE92AFFFFFFFFFFFFFFFFFFF969FFFFFFFFFFFFFAABFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_0C = 256'hFFFFFF9AFFFFFFFFFFFFFC0014047FFFFFFFFFFFFFFFFFF96A54D5F5C6ABFFFF;
defparam sdpb_inst_10.INIT_RAM_0D = 256'h9A6925BDE16ABFFFFFFFFFFFF82BFFFA86BFFFFFFFFFFFFFFFFFFFE555FFFFFF;
defparam sdpb_inst_10.INIT_RAM_0E = 256'hFFFFFFFF91AFFFFFFFFFFFEAAFFFFFFFFFFFFFF0E80100FFFFFFFFFFFFFFFFFE;
defparam sdpb_inst_10.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFE96AA546D1716AAFFFFFFFFFFFE56FFFE9DBFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_10 = 256'hA96AFFFFFFFFFFFFFFFFFFFFFE555FFFFFFFFFFAAAFFFFFFFFFFFFFFC002408F;
defparam sdpb_inst_10.INIT_RAM_11 = 256'hFFFFFFFFFF0F80001FFFFFFFFFFFFFFF96A655A6CA716AAFFFFFFFFFFFA0AFFF;
defparam sdpb_inst_10.INIT_RAM_12 = 256'hBFFFFFFFFFF95AFFFA46AFFFFFFFFFFFFFFFFFFFFFF9166FFFFFFFE6AABFFFFF;
defparam sdpb_inst_10.INIT_RAM_13 = 256'h55BBFF5599AFFFFFFFFFFFFFFFBC0034083FFFFFFFFFFFFFEAAA55D97DAA85AA;
defparam sdpb_inst_10.INIT_RAM_14 = 256'hFA6A97E9E46AA416ABFFFFFFFFFF82BFFEA5AAFFFFFFFFFFFFFFFFFFFFFFE855;
defparam sdpb_inst_10.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFA444555556556BFFFFFFFFFFFFFFFEF0B80100FFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_16 = 256'h3040C3FFFFFFFFFFFEBAA5BD5EB6AA986ABFFFFFFFFFE56FFEA85ABFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_17 = 256'hFFEA96AAFFFFFFFFFFFFFFFFFFFADBFEA0341555546FFFFFFFFFFFFFFFFFFBC0;
defparam sdpb_inst_10.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFEF0B80000FFFFFFFFFFFE96979555B5AA9B5ABFFFFFFFFFAFB;
defparam sdpb_inst_10.INIT_RAM_19 = 256'h9B5ABFFFFFFFFFA1BFFAA86AAFFFFFFFFFFFFFEFEAAA93A9ABAA545151AFFFFF;
defparam sdpb_inst_10.INIT_RAM_1A = 256'hAA7BEAAAAAFFFFFFFFFFFFFFFFFFFFFFBC030000FFFFFFFFFFEA95571555B6AA;
defparam sdpb_inst_10.INIT_RAM_1B = 256'hFFFEA555F155EBAAA8B2ABFFFFFFFFF86BFEAA5AABFFFFFFFFFFFFFAEAAA876A;
defparam sdpb_inst_10.INIT_RAM_1C = 256'hFFFFFBEAAAAA98AAAAAA7ABEBFFFFFFFFFFFFFFFFFFFFFFFFEF0B8000FFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1D = 256'hFFFBC00000BFFFFFFFFFA9E657DAABDAAA576AABFFFFFFFE82BAAAA5AAAAFFFF;
defparam sdpb_inst_10.INIT_RAM_1E = 256'hE86FEAA95AAAEFFFBFFFFABAAAAA969ABAAAAB4ABFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFEF00000FFFFFFFFFF9E2556F28B6AA9986AAFFFFFFFB;
defparam sdpb_inst_10.INIT_RAM_20 = 256'hAAB251AAAFFFFFFFFE4AAAAA96AAABFFFFFFFFEAAAAA9596AFAAAAA7AAFFFFFF;
defparam sdpb_inst_10.INIT_RAM_21 = 256'hBBFEAAAA96AAFFFFFFFFFFFFFFFFFFFFFFFFFFDC0002FFFFFFFFF600D6693FFD;
defparam sdpb_inst_10.INIT_RAM_22 = 256'hFFFFF9829D96A969AAA4576AAAFFFFFFFFA1AAAAA96AAABBFFFFBFFEAAAAA565;
defparam sdpb_inst_10.INIT_RAM_23 = 256'hFFFFFFFEEAAAA95B7FFFF8AFAA9EEBFFFFFFFFFFFFFFFFFFFFFFFFFF8502BFFF;
defparam sdpb_inst_10.INIT_RAM_24 = 256'hFFFFFFFFFFEABFFFFFFFF86053D6AAA96AA915C6AABFBFFFFFFA0AAAAA96AABE;
defparam sdpb_inst_10.INIT_RAM_25 = 256'hFFFFA1AAAAA96AABAFBFFFFAFAAAAA545BFFFC58FFA9CE7BFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_26 = 256'hBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA5656A19AAAAAAA7775AAABEFFF;
defparam sdpb_inst_10.INIT_RAM_27 = 256'h656A912C6AAAFBFFFAFBA92AAAAA96AAAAFFBFEAEAAAAA952DBFFFD5583CAD8E;
defparam sdpb_inst_10.INIT_RAM_28 = 256'h496EFFF55158FC95CEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE95655A5669;
defparam sdpb_inst_10.INIT_RAM_29 = 256'hFFFFFEA55595AD565C55A9E71AAAAAEBFFEBEA89AAAAA76AAAABAEEAAAAAAAA5;
defparam sdpb_inst_10.INIT_RAM_2A = 256'hAAAAAABAAAAAAAA9509BBFFC545519FA97F7BFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFAA555A556D69E6569EB5AAAAABFFEFFEA9EAAAAA56;
defparam sdpb_inst_10.INIT_RAM_2C = 256'hAAAFABAA82AAAAA56AAAAAAAAAAAAAAA942E7FFFD5555559EAEFD9BFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_2D = 256'h5AFA2ABABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEA69765656996A69D9E85AAAAA;
defparam sdpb_inst_10.INIT_RAM_2E = 256'hAABEA6A15E85AAAAAAAAAAAAA86AAAAA5AAAAAAAAAAAAAAAA544BF7FF5515455;
defparam sdpb_inst_10.INIT_RAM_2F = 256'hAA53BEFFBD545515456EFAA0BAFFFFFFFFFFFFFFFFFFFFFFFFFFEEFAA569D5C0;
defparam sdpb_inst_10.INIT_RAM_30 = 256'hFFFFFFAAA8559540002B5AAA95EC6AAAAAAAAAAAAA46AAAAA9AAAAAAAAAAAAAA;
defparam sdpb_inst_10.INIT_RAM_31 = 256'hAB1AAAAAAAAAAAAAAA9517FFFF155555515BFFFAC6A2FFFFFFFFFFFFFFFFFFFF;
defparam sdpb_inst_10.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFBEA95559400000A5AA95BC6AAAAAAAAAAAAA56AAA;
defparam sdpb_inst_10.INIT_RAM_33 = 256'hAAAAAAAAAAAAF6AAAA95AAAAAAAAAAAAAAA951FBF0CFD5555555FFBFFFC62AFF;
defparam sdpb_inst_10.INIT_RAM_34 = 256'h1545700FFFFFC2AA8BAAFFFFFFFFFFFEFFFFFFFEEAA9556AAAAAC56AAAA54C6A;
defparam sdpb_inst_10.INIT_RAM_35 = 256'hAAAAAAB2AAAA85C6AAAAAAAAAAAAAD6AAAA55AAAAAAAAAAAAAAA94E7BF0E23C5;
defparam sdpb_inst_10.INIT_RAM_36 = 256'hAAAAA94E56FFB333D1515C030F3FFF49A52AFFFFFFFFFFFFFFFFFFFBFEAAB55A;
defparam sdpb_inst_10.INIT_RAM_37 = 256'hFFFFFFFFAEEAA9559AAAAAAAAAAAAB6DAAAAAAAAAAAAAA16AAAA76AAAAAAAAAA;
defparam sdpb_inst_10.INIT_RAM_38 = 256'h6AAA946AAAAAAAAAAAAAAA94E95AEAAC3C2555008000FFFCC45AAAAAEFFFEFFF;
defparam sdpb_inst_10.INIT_RAM_39 = 256'h9529BAAAAEFFFBBFFFFFFFFBEBFAAAA15AAAAAAAAAAAAA6A1AAAAAAAAAAAAA91;
defparam sdpb_inst_10.INIT_RAM_3A = 256'h71AAAAAAAAAAAAA996AAA956AAAAAAAAAAAAAAA953956FEAAB3C3570000000CF;
defparam sdpb_inst_10.INIT_RAM_3B = 256'hEAAAFC3000000000F54158AAAAAAFFFAFFBFEFEBFAAAAAAA456AAAAAAAAAABD5;
defparam sdpb_inst_10.INIT_RAM_3C = 256'hA915AAAAAAAAAAA1786AAAAAAAAAAAAAB56AAA8D6AAAAAAAAAAAAAAA9539556B;
defparam sdpb_inst_10.INIT_RAM_3D = 256'hAAAAAAAAA954E5998ECEAAF83CC000000F6551559AAAAEFFFAFEFFFBBBEBAAAA;
defparam sdpb_inst_10.INIT_RAM_3E = 256'hAABEFEEEAAAEAEAAAA9656BAAAAAAAF056D6AAAAAAAAAAAAA856AAA516AAAAAA;
defparam sdpb_inst_10.INIT_RAM_3F = 256'hAA416AAA55AAAAAAAAAAAAAAAAA543931EBE3ED0FB30000000C69AA56FAAAAAA;

SDPB sdpb_inst_11 (
    .DO({sdpb_inst_11_dout_w[29:0],sdpb_inst_11_dout[7:6]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[14],ada[13]}),
    .BLKSELB({gw_gnd,adb[14],adb[13]}),
    .ADA({ada[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]}),
    .ADB({adb[12:0],gw_gnd})
);

defparam sdpb_inst_11.READ_MODE = 1'b1;
defparam sdpb_inst_11.BIT_WIDTH_0 = 2;
defparam sdpb_inst_11.BIT_WIDTH_1 = 2;
defparam sdpb_inst_11.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_11.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_11.RESET_MODE = "SYNC";
defparam sdpb_inst_11.INIT_RAM_00 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAA55511456AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_01 = 256'hAAAAAAAAAAAAAAAA80116AAAAAAAAAAAAAAAA6AAAAAA2AAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_02 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95154155AAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_03 = 256'h11456AAAAAAAAAAAAAAAAAAAAAAAAAAAA0001AAAAAAAAAAAAAAAA9AAAAAA8AAA;
defparam sdpb_inst_11.INIT_RAM_04 = 256'hAAAAAA9AAAAAA2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA554;
defparam sdpb_inst_11.INIT_RAM_05 = 256'hAAAAAAAAAAAAAA95154151AAAAAAAAAAAAAAAAAAAAAAAAAAA91005AAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_06 = 256'hAA80116AAAAAAAAAAAAAAAA6AAAAA86AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_07 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55411456AAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_08 = 256'hAAAAAAAAAAAAAAAAAAA0041AAAAAAAAAAAAAAAA9AAAAAA5AAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_09 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA95554151AAAAAAA;
defparam sdpb_inst_11.INIT_RAM_0A = 256'hAAA45415456AAAAAAAAAAAAAAAAAAAAAAAA80005AAAAAAAAAAAAAAAA5AAAAAA2;
defparam sdpb_inst_11.INIT_RAM_0B = 256'hAAAAAAAAA6AAAAA8AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_0C = 256'hAAAAAAAAAAAAAAAAAAAA91554151AAAAAAAAAAAAAAAAAAA9555600016AAAAAAA;
defparam sdpb_inst_11.INIT_RAM_0D = 256'h555540001AAAAAAAAAAAAAAAA9AAAAAA2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_0E = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA45015456AAAAAAAAAAAAAAAAA9;
defparam sdpb_inst_11.INIT_RAM_0F = 256'hAAAAAAAAAAAAAAAA5555510045AAAAAAAAAAAAAAAA9AAAAAA2AAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_10 = 256'hA8AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA915541516;
defparam sdpb_inst_11.INIT_RAM_11 = 256'hAAAAAAAAA45015455AAAAAAAAAAAAAAA95555400155AAAAAAAAAAAAAAAA6AAAA;
defparam sdpb_inst_11.INIT_RAM_12 = 256'hAAAAAAAAAAAA6AAAAA6AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_13 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAA915541516AAAAAAAAAAAAAA555550001556AAA;
defparam sdpb_inst_11.INIT_RAM_14 = 256'hAA555400015555AAAAAAAAAAAAAA9AAAAAA2AAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_15 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA45015455AAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_16 = 256'h451516AAAAAAAAAAAA95550000055556AAAAAAAAAAAAA9AAAAA9AAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_17 = 256'hAAAA8AAAAAAAAAAAAAAAAAAAAAAA95AAAA9AAAAAAAAAAAAAAAAAAAAAAAAAA915;
defparam sdpb_inst_11.INIT_RAM_18 = 256'hAAAAAAAAAAAAAAA45015456AAAAAAAAAAAA95540000055551AAAAAAAAAAAAA1A;
defparam sdpb_inst_11.INIT_RAM_19 = 256'h51AAAAAAAAAAAAA6AAAAA6AAAAAAAAAAAAAAAAAAAAAAA4556AAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_1A = 256'h555AAAAAAAAAAAAAAAAAAAAAAAAAAAAA91545155AAAAAAAAAAAA955440000555;
defparam sdpb_inst_11.INIT_RAM_1B = 256'hAAAAA51504000055551AAAAAAAAAAAAA6AAAAA2AAAAAAAAAAAAAAAAAAAAAA455;
defparam sdpb_inst_11.INIT_RAM_1C = 256'hAAAAAAAAAAAAA51555555AAAAAAAAAAAAAAAAAAAAAAAAAAAAA4501555AAAAAAA;
defparam sdpb_inst_11.INIT_RAM_1D = 256'hAAA9155555AAAAAAAAAAA954540000155545AAAAAAAAAAAA9AAAAAA2AAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_1E = 256'hA9AAAAAA6AAAAAAAAAAAAAAAAAAAA9155555556AAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_1F = 256'hAAAAAAAAAAAAAAAAAAAAA455555AAAAAAAAAA9595540410555506AAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_20 = 256'h55541AAAAAAAAAAAAA9AAAAA9AAAAAAAAAAAAAAAAAAAAA45555555556AAAAAAA;
defparam sdpb_inst_11.INIT_RAM_21 = 256'h55555555556AAAAAAAAAAAAAAAAAAAAAAAAAAAA15556AAAAAAAAA9AA55554001;
defparam sdpb_inst_11.INIT_RAM_22 = 256'hAAAAA96955555555555505AAAAAAAAAAAAA9AAAAA8AAAAAAAAAAAAAAAAAAAA91;
defparam sdpb_inst_11.INIT_RAM_23 = 256'hAAAAAAAAAAAAAAA45555515555556AAAAAAAAAAAAAAAAAAAAAAAAAAAA555AAAA;
defparam sdpb_inst_11.INIT_RAM_24 = 256'hAAAAAAAAAAAAAAAAAAAAA95A545555555555416AAAAAAAAAAAAA6AAAAA8AAAAA;
defparam sdpb_inst_11.INIT_RAM_25 = 256'hAAAAA6AAAAA8AAAAAAAAAAAAAAAAAAAA55555501555515AAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_26 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA55540555555555405AAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_27 = 256'h55555456AAAAAAAAAAAAAA6AAAAA8AAAAAAAAAAAAAAAAAAA9155554001965015;
defparam sdpb_inst_11.INIT_RAM_28 = 256'hA45555500001564015AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9555005555;
defparam sdpb_inst_11.INIT_RAM_29 = 256'hAAAAAAA55500015551555505AAAAAAAAAAAAAAA6AAAAA8AAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_2A = 256'hAAAAAAAAAAAAAAAAA9555554000001550005AAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_2B = 256'hAAAAAAAAAAAAAAAAAAAAAAA855400001550055505AAAAAAAAAAAAAA96AAAAA6A;
defparam sdpb_inst_11.INIT_RAM_2C = 256'hAAAAAAAA9AAAAAA2AAAAAAAAAAAAAAAAAA90555500000001550006AAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_2D = 256'h01554016AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA414050001140001506AAAAAA;
defparam sdpb_inst_11.INIT_RAM_2E = 256'h00000005506AAAAAAAAAAAAAA9AAAAAA2AAAAAAAAAAAAAAAAAA1055550000000;
defparam sdpb_inst_11.INIT_RAM_2F = 256'hAAA94155540000000015550516AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA0001515;
defparam sdpb_inst_11.INIT_RAM_30 = 256'hAAAAAAAAAA001555554000001506AAAAAAAAAAAAAA9AAAAAA2AAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_31 = 256'hA8AAAAAAAAAAAAAAAAAA94155540000000015555141AAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_32 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAA9000155555500001506AAAAAAAAAAAAAA9AAAA;
defparam sdpb_inst_11.INIT_RAM_33 = 256'hAAAAAAAAAAAA5AAAAA8AAAAAAAAAAAAAAAAAA8055A6540000000555555145AAA;
defparam sdpb_inst_11.INIT_RAM_34 = 256'h00001AA55555145AAAAAAAAAAAAAAAAAAAAAAAAAAAA9000000001540000516AA;
defparam sdpb_inst_11.INIT_RAM_35 = 256'h000000040000116AAAAAAAAAAAAAA2AAAAA8AAAAAAAAAAAAAAAAAA5455A59950;
defparam sdpb_inst_11.INIT_RAM_36 = 256'hAAAAAAA555555999500002A9A595555058AAAAAAAAAAAAAAAAAAAAAAAAAA9000;
defparam sdpb_inst_11.INIT_RAM_37 = 256'hAAAAAAAAAAAAAA000000000000000016AAAAAAAAAAAAAA6AAAAA5AAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_38 = 256'hAAAAA2AAAAAAAAAAAAAAAAAA55555556969000AA6AAA5555500AAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_39 = 256'h40501AAAAAAAAAAAAAAAAAAAAAAAAAA40000000000000001AAAAAAAAAAAAAAA6;
defparam sdpb_inst_11.INIT_RAM_3A = 256'h5AAAAAAAAAAAAAAA6AAAAA2AAAAAAAAAAAAAAAAAA95555555596901AAAAAAA65;
defparam sdpb_inst_11.INIT_RAM_3B = 256'h55555696AAAAAAAA5000155AAAAAAAAAAAAAAAAAAAAAAAAA9000000000000100;
defparam sdpb_inst_11.INIT_RAM_3C = 256'hAA4000000000004406AAAAAAAAAAAAAA8AAAAA96AAAAAAAAAAAAAAAAAA955555;
defparam sdpb_inst_11.INIT_RAM_3D = 256'hAAAAAAAAAAAA541565655556966AAAAAA50000055AAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_3E = 256'hAAAAAAAAAAAAAAAAAAA9001000000014016AAAAAAAAAAAAAA9AAAAA8AAAAAAAA;
defparam sdpb_inst_11.INIT_RAM_3F = 256'hAA9AAAAA8AAAAAAAAAAAAAAAAAAAA95015559500559AAAAAAA500000155AAAAA;

SDPB sdpb_inst_12 (
    .DO({sdpb_inst_12_dout_w[27:0],sdpb_inst_12_dout[3:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_12.READ_MODE = 1'b1;
defparam sdpb_inst_12.BIT_WIDTH_0 = 4;
defparam sdpb_inst_12.BIT_WIDTH_1 = 4;
defparam sdpb_inst_12.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_12.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_12.RESET_MODE = "SYNC";
defparam sdpb_inst_12.INIT_RAM_00 = 256'hBDCA9751C6CD18B983CA48724794AE23D398AC1C1568AA9AAABBAAAAA9998997;
defparam sdpb_inst_12.INIT_RAM_01 = 256'h865340A802459AB71547F4107BCADDCF0EFEEFFECEEE0EFEEFEFFFFEDDFDFDFD;
defparam sdpb_inst_12.INIT_RAM_02 = 256'h99AA99998A988988877665421DA4C065C65C1DDBB01BADE0EC0BC83188778996;
defparam sdpb_inst_12.INIT_RAM_03 = 256'h5B06A3B1B0568989A9A9AA989999988777543B73E7D112421CD26E2257889989;
defparam sdpb_inst_12.INIT_RAM_04 = 256'hCDCDDDEEEEDEEEE0DDF0EFEEFEFFECFCEEB99AA8642D8265279182A1AEDE72DE;
defparam sdpb_inst_12.INIT_RAM_05 = 256'h5A16FF7B98F77A99EE0FCA01D731898B9A86521EF71359E0EB5C56F02FB789BC;
defparam sdpb_inst_12.INIT_RAM_06 = 256'h766441DEF202AE3210EB4A8F34575887788889999899A998887887666420D82C;
defparam sdpb_inst_12.INIT_RAM_07 = 256'hDEDCCCBBAA8743EA70AB808BC0C5CF61EE6D97E12CF35898989A9A9999898878;
defparam sdpb_inst_12.INIT_RAM_08 = 256'hA99984010A9E288CEFEB57FAA101FED6DBECCDDEEEDDDADEEEDC0EED0DFEFFDE;
defparam sdpb_inst_12.INIT_RAM_09 = 256'h7877799898998988878867667654310B84EA1761AD6E88F3E89B085A6D9C5E08;
defparam sdpb_inst_12.INIT_RAM_0A = 256'h8E6CC2CEB6D1448889988989898888777857642EBB08BE8DF0FE5E3D9E245887;
defparam sdpb_inst_12.INIT_RAM_0B = 256'h3A88BCDDDCEEDECBDEDEBEEEECDCDEFCCDBCCCABEBAB977642FC5D9DE6D7FE3C;
defparam sdpb_inst_12.INIT_RAM_0C = 256'h1FCA61D6D2214D98BAF33F2F8462459DC1B68A6610EFE016BBFCB92AFFB1021D;
defparam sdpb_inst_12.INIT_RAM_0D = 256'h865656300C5BFEF09CFED89140BF245676777788897989998878877676764441;
defparam sdpb_inst_12.INIT_RAM_0E = 256'hCDDCCDBEDCCAABB9876330EB83E70594A2270F94E5AF23577998788988888877;
defparam sdpb_inst_12.INIT_RAM_0F = 256'hAACCEFD6500CE78E29CEEAA4BE61D1000C3D68AABDCCCDDCCCBCCCDBCCCCCBCC;
defparam sdpb_inst_12.INIT_RAM_10 = 256'h667677778786777887777777767656555320DFB751A49DE6BBFDEC1D934B5089;
defparam sdpb_inst_12.INIT_RAM_11 = 256'hE9A86BD069BF134577779979787778777767555332FBB537439ECB7B00FEA023;
defparam sdpb_inst_12.INIT_RAM_12 = 256'h020C38269ABCBCBCDDCBBCBCBBBCDBACDABCDABACCCCAB9AA997876342FDA64F;
defparam sdpb_inst_12.INIT_RAM_13 = 256'h56433201DC9840807BF357CDFEEA532B97712030BDEFBB6A5F5CEDBB527E32F1;
defparam sdpb_inst_12.INIT_RAM_14 = 256'h77666654432FDA714EC5BAB823E470AF24686778777777877878678667677766;
defparam sdpb_inst_12.INIT_RAM_15 = 256'hABBCADBAAC9DCC9AA9AAA9876655420FDCCA9AACDEFF24457667787887977858;
defparam sdpb_inst_12.INIT_RAM_16 = 256'hE57DDEE0E5163AA74A7C2ACBB828DF36323F2D5A9C79ABAACCDBDCBCDCBBCBBA;
defparam sdpb_inst_12.INIT_RAM_17 = 256'hB045566667665778666577765766766675655443210ECB86209057CFFB1D0FD0;
defparam sdpb_inst_12.INIT_RAM_18 = 256'h4321111F0011334568777777776776776677656654421EC89FC709CCC926DEF2;
defparam sdpb_inst_12.INIT_RAM_19 = 256'h5DE23F0451A4D6A89AABBBBA9ACADBBBBACABAAA9A9ABACAA9A9A99988787754;
defparam sdpb_inst_12.INIT_RAM_1A = 256'h5555654443000FFECA862FB1469ABC113EE1381CF0FF0D9B49A77B428AA607F2;
defparam sdpb_inst_12.INIT_RAM_1B = 256'h6574555655454320EA2A5D7CFDB8FBD657D13446655557667566766656555656;
defparam sdpb_inst_12.INIT_RAM_1C = 256'hCAAABAAABAA9BB9B9AA9A9A99989898976656444513344545656777775666676;
defparam sdpb_inst_12.INIT_RAM_1D = 256'h134441C46E20122F2FD36760165B95D292FD2342219CE9D599999CAB9C8BBCAC;
defparam sdpb_inst_12.INIT_RAM_1E = 256'hEEC8F144446557566565665766564555664545565544323100FDCA9643803784;
defparam sdpb_inst_12.INIT_RAM_1F = 256'h97775666454443456556566756665466666666555442553310EDA89BEDFEC6C0;
defparam sdpb_inst_12.INIT_RAM_20 = 256'hD2453235333109D02379999A9AAA8AABBA9999AA999BA8999999998987799887;
defparam sdpb_inst_12.INIT_RAM_21 = 256'h45555655555444231321F0FDDCB861B38C66848530C40BDFEF0DF14540367996;
defparam sdpb_inst_12.INIT_RAM_22 = 256'h455455544444452332232FFDEF000EC53EF71BF2345465455454554544655555;
defparam sdpb_inst_12.INIT_RAM_23 = 256'hAABAA989899AAA99999A99977878789978887767566656565564556567566754;
defparam sdpb_inst_12.INIT_RAM_24 = 256'h73F9E19D834441B8B9D314A3716BE46A833D3B425454320AB50078AAAAB997A9;
defparam sdpb_inst_12.INIT_RAM_25 = 256'hE99D5D9F033423455544544544453354434545555554455443343010F0DFECB8;
defparam sdpb_inst_12.INIT_RAM_26 = 256'h6778777776666566555564655576445445454433444444423333321110000FE1;
defparam sdpb_inst_12.INIT_RAM_27 = 256'h5861401C446453322DB7F16677A8999AB999998A978888898988788768777777;
defparam sdpb_inst_12.INIT_RAM_28 = 256'h432343445544444444443333212220F0FDCB750A2C6A95543FABFA14E40B28BC;
defparam sdpb_inst_12.INIT_RAM_29 = 256'h3434333433323333223323110110111011FDB16CF12133344234513434433444;
defparam sdpb_inst_12.INIT_RAM_2A = 256'h988898A889888877778777867776676777777767656757766675557655646453;
defparam sdpb_inst_12.INIT_RAM_2B = 256'h12200EEB862C0A59A2552FC93DCCDCA3BC15164296566456311EA5E255788798;
defparam sdpb_inst_12.INIT_RAM_2C = 256'h211100FFF0F13313223222123434244223233344432433433334543333324443;
defparam sdpb_inst_12.INIT_RAM_2D = 256'h656666767576667555544556644754534354233343123121231214321F011012;
defparam sdpb_inst_12.INIT_RAM_2E = 256'h2E4C89A32A95565354322EB9F146677777897899999877676786866657777556;
defparam sdpb_inst_12.INIT_RAM_2F = 256'h12222232213223233433432322324334333332200FDB8418E53792532E250C5C;
defparam sdpb_inst_12.INIT_RAM_30 = 256'h433333223112F120122212222111221110101101000102111213112222323234;
defparam sdpb_inst_12.INIT_RAM_31 = 256'h5868885877787768867687673566658645454675566555556544555556455454;
defparam sdpb_inst_12.INIT_RAM_32 = 256'h3444343331210FFB94059163D3330308540A134218572356421222E853004667;
defparam sdpb_inst_12.INIT_RAM_33 = 256'h0110F1F01011111F0123FF02120322F1112011320F1231331321222233322222;
defparam sdpb_inst_12.INIT_RAM_34 = 256'h4554443655553564444558342433444435124212213F33001210112011310101;
defparam sdpb_inst_12.INIT_RAM_35 = 256'h54C100AFC6E6255654534318F70CF23467867777677888687567666686774564;
defparam sdpb_inst_12.INIT_RAM_36 = 256'h120111110111F01111103222222222333333444335343322F0DB73D46F51B42F;
defparam sdpb_inst_12.INIT_RAM_37 = 256'h44342211101012010010FFF102F111F00000100011000111110210111111F200;
defparam sdpb_inst_12.INIT_RAM_38 = 256'h3446666866668766877656556656254445544445245433554544534335344542;
defparam sdpb_inst_12.INIT_RAM_39 = 256'h22334443445455434311FCCA61A23D813510C9F4ABEA65353465432330F7EB03;
defparam sdpb_inst_12.INIT_RAM_3A = 256'h0F0F000FFFFF0F0F01FFFF100001F111000FF0F0F0FFFFF01F00011101110221;
defparam sdpb_inst_12.INIT_RAM_3B = 256'h443344323343234342443433333233343334322110000FF0FFFE1FFEFF0F01FF;
defparam sdpb_inst_12.INIT_RAM_3C = 256'h1E89C5E65FA0F9744555574121F0DEAC12365557666557576663555654676654;
defparam sdpb_inst_12.INIT_RAM_3D = 256'hFFFFFFFF0EFE0FF0EF0FEEE0000111101122222444556446644434110EC74F8F;
defparam sdpb_inst_12.INIT_RAM_3E = 256'h2332231211000FEFFEFFFEFFEEFFFF0FFFF0E0FFFFFEE1E00FE0EFFF00FFFFFF;
defparam sdpb_inst_12.INIT_RAM_3F = 256'hBF12444655666556566554665443344422333322325222233223223333323133;

SDPB sdpb_inst_13 (
    .DO({sdpb_inst_13_dout_w[27:0],sdpb_inst_13_dout[7:4]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd})
);

defparam sdpb_inst_13.READ_MODE = 1'b1;
defparam sdpb_inst_13.BIT_WIDTH_0 = 4;
defparam sdpb_inst_13.BIT_WIDTH_1 = 4;
defparam sdpb_inst_13.BLK_SEL_0 = 3'b110;
defparam sdpb_inst_13.BLK_SEL_1 = 3'b110;
defparam sdpb_inst_13.RESET_MODE = "SYNC";
defparam sdpb_inst_13.INIT_RAM_00 = 256'hAAAAAAAA99841112747732272235452101115799AAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_01 = 256'h8888887133333333321167765AAAAAAABAAAAAAAAAAABAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_02 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAA999887634516575576200010010677888888888;
defparam sdpb_inst_13.INIT_RAM_03 = 256'h102126799AAAAAAAAAAAAAAAAAAAAAAAAAAAA911899AAAAAA91899AAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_04 = 256'hAAAAAAAAAAAAAAABAAABAAAAAAAAAAAAAAAAAAAAAAA999842112232366626410;
defparam sdpb_inst_13.INIT_RAM_05 = 256'h877503505566566300100012675888888888888721333334333210677665AAAA;
defparam sdpb_inst_13.INIT_RAM_06 = 256'hAAAAAA96018999AAAA991899AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9998;
defparam sdpb_inst_13.INIT_RAM_07 = 256'hAAAAAAAAAAAAAA99998642111212222110211568999AAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_08 = 256'h8888888887123333333332007777665AAAAAAAAAAAAAAAAAAAAABAAABAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_09 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA999888765006355565742111211102768;
defparam sdpb_inst_13.INIT_RAM_0A = 256'h13211567899AAAAAAAAAAAAAAAAAAAAAAAAAAAA9911178999A99917899AAAAAA;
defparam sdpb_inst_13.INIT_RAM_0B = 256'h45AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99988754444210;
defparam sdpb_inst_13.INIT_RAM_0C = 256'hA999998877654355555667401111110028688888887113333333333100677776;
defparam sdpb_inst_13.INIT_RAM_0D = 256'hAAAAAAAAA9900679999999217999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_0E = 256'hAAAAAAAAAAAAAAAAAAAAAA9999888765334566788999AAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_0F = 256'h1110567888871122333333332011577776437AAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_10 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9999998876554545556567411310;
defparam sdpb_inst_13.INIT_RAM_11 = 256'h888888899999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9971178999999811689AAA;
defparam sdpb_inst_13.INIT_RAM_12 = 256'h7776474AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA999998;
defparam sdpb_inst_13.INIT_RAM_13 = 256'hAAAAAAAA99999988765535455555762200111121767772122233333333101147;
defparam sdpb_inst_13.INIT_RAM_14 = 256'hAAAAAAAAAAA999111789999998017999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_15 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9999999999999AAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_16 = 256'h710100010116673122223333333200107766763774AAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_17 = 256'h9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA999999988765355556556;
defparam sdpb_inst_13.INIT_RAM_18 = 256'hAAAAAAA9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9991068999999970279;
defparam sdpb_inst_13.INIT_RAM_19 = 256'h1167767648776AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_1A = 256'hAAAAAAAAAAAAA999999998887655555665568610010011531122223333333101;
defparam sdpb_inst_13.INIT_RAM_1B = 256'hAAAAAAAAAAAAAAAA9998889999998504899AAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_1C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_1D = 256'h54666656871111102401222333333321010677777763175AAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_1E = 256'h06899AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99999999887655;
defparam sdpb_inst_13.INIT_RAM_1F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99999999999981;
defparam sdpb_inst_13.INIT_RAM_20 = 256'h21111777777776666AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_21 = 256'hAAAAAAAAAAAAAAAAAAAA9A999999998876554466665685000011611223333333;
defparam sdpb_inst_13.INIT_RAM_22 = 256'hAAAAAAAAAAAAAAAAAAAAA99999AAA9998007999AAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_23 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_24 = 256'h998877554466665672011137112223333320107777777776666AAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_25 = 256'h99833899AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9A999999;
defparam sdpb_inst_13.INIT_RAM_26 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99A;
defparam sdpb_inst_13.INIT_RAM_27 = 256'h333311137777777776665AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_28 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9A99999998865545666556711101701222;
defparam sdpb_inst_13.INIT_RAM_29 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9999999AAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_2A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_2B = 256'hAAAAA99999988655466665567001060122333211077777777776675AAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_2C = 256'hAAAAAA999A9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_2D = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAA;
defparam sdpb_inst_13.INIT_RAM_2E = 256'h5012221110777777777776668AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_2F = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99999987655466665564010;
defparam sdpb_inst_13.INIT_RAM_30 = 256'hAAAAAAAAAAAA9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_31 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_32 = 256'hAAAAAAAAAAAAA999999876554666651111121111103767777777775666AAAAAA;
defparam sdpb_inst_13.INIT_RAM_33 = 256'hAAAA9A9AAAAAAAA9AAAA99AAAAAAAA9AAAAAAAAAA9AAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_34 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_35 = 256'h41451500004777767777777626769AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_36 = 256'hAAAAAAAAAAAA9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9A99998875555665;
defparam sdpb_inst_13.INIT_RAM_37 = 256'hAAAAAAAAAAAAAAAAAAAA999AAA9AAA9AAAAAAAAAAAAAAAAAAAAAAAAAAAAA9AAA;
defparam sdpb_inst_13.INIT_RAM_38 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_39 = 256'hAAAAAAAAAAAAAAAAAAAA999999887555666655565777777777677777776659AA;
defparam sdpb_inst_13.INIT_RAM_3A = 256'hA9A9AAA99999A9A9AA9999AAAAAA9AAAAAA99A9A9A99999AA9AAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_3B = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99A9999A99999A9AA99;
defparam sdpb_inst_13.INIT_RAM_3C = 256'h75555655546877777777767777676659AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam sdpb_inst_13.INIT_RAM_3D = 256'h99999999A999A99A99A9999AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9999887;
defparam sdpb_inst_13.INIT_RAM_3E = 256'hAAAAAAAAAAAAA99999999999999999A9999A9A9999999A9AA99A9999AA999999;
defparam sdpb_inst_13.INIT_RAM_3F = 256'h99AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;

SDPB sdpb_inst_14 (
    .DO({sdpb_inst_14_dout_w[23:0],sdpb_inst_14_dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,lut_f_0}),
    .BLKSELB({gw_gnd,gw_gnd,lut_f_1}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_14.READ_MODE = 1'b1;
defparam sdpb_inst_14.BIT_WIDTH_0 = 8;
defparam sdpb_inst_14.BIT_WIDTH_1 = 8;
defparam sdpb_inst_14.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_14.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_14.RESET_MODE = "SYNC";
defparam sdpb_inst_14.INIT_RAM_00 = 256'h938E867B716351561E13655456577179757474747674736F6B73727170706959;
defparam sdpb_inst_14.INIT_RAM_01 = 256'h9FA1A0A1A1A1A2A2A2A2A3A4A4A5A4A4A4A5A4A5A5A4A4A4A3A3A2A19F9E9A97;
defparam sdpb_inst_14.INIT_RAM_02 = 256'h9E9F9F9F9E9F9F9E9E9E9E9E9E9E9E9E9E9E9E9E9F9E9E9E9EA09F9F9FA09FA0;
defparam sdpb_inst_14.INIT_RAM_03 = 256'h9D9E9C9F9E9E9E9E9E9E9E9F9D9F9EA09E9F9F9E9F9F9E9F9F9E9E9E9F9F9F9D;
defparam sdpb_inst_14.INIT_RAM_04 = 256'hA2A2A2A2A3A1A2A2A2A09F9F9F9F9F9C9E9F9EA09D9F9F9E9D9E9D9D9D9D9E9E;
defparam sdpb_inst_14.INIT_RAM_05 = 256'hA3A1A2A1A1A1A3A2A2A1A1A1A1A1A3A1A0A2A1A2A1A2A2A1A2A2A3A4A3A0A2A1;
defparam sdpb_inst_14.INIT_RAM_06 = 256'h647F9AA0A1A2A4A4A4A5A5A5A4A5A4A5A5A4A5A5A5A5A5A5A4A4A3A4A4A3A3A2;
defparam sdpb_inst_14.INIT_RAM_07 = 256'h9E9C9A96908B827870664C1128120B58585C7073757274715550856C70706D64;
defparam sdpb_inst_14.INIT_RAM_08 = 256'h9F9F9FA09FA0A1A0A1A1A2A1A3A4A2A4A5A4A6A4A4A5A6A6A6A6A5A5A4A4A2A1;
defparam sdpb_inst_14.INIT_RAM_09 = 256'h9E9C9E9E9C9D9F9D9F9D9E9E9D9D9D9D9E9D9C9D9E9D9D9D9D9D9E9E9F9F9E9E;
defparam sdpb_inst_14.INIT_RAM_0A = 256'h9E9C9C9C9E9E9D9E9F9F9D9D9D9D9E9F9D9E9D9D9E9F9D9D9D9D9D9E9E9D9E9E;
defparam sdpb_inst_14.INIT_RAM_0B = 256'hA1A0A1A1A1A1A2A2A0A0A1A09E9D9E9E9E9D9D9D9D9D9D9D9C9C9D9D9D9C9C9C;
defparam sdpb_inst_14.INIT_RAM_0C = 256'hA2A2A0A1A2A1A1A2A0A2A1A0A1A0A0A0A1A2A1A2A0A1A0A1A2A0A2A1A0A1A09F;
defparam sdpb_inst_14.INIT_RAM_0D = 256'h6B695B9D9DA0A1A3A4A5A4A5A5A4A4A5A3A4A4A3A4A4A4A5A5A5A3A4A4A3A4A3;
defparam sdpb_inst_14.INIT_RAM_0E = 256'hA4A2A0A09E9B99968D8A817C756756693D13735D60636F736D2F737E7E736C6E;
defparam sdpb_inst_14.INIT_RAM_0F = 256'h9C9D9F9FA09E9F9EA0A0A0A1A3A2A2A3A4A4A4A4A5A3A5A6A5A6A6A6A6A6A5A5;
defparam sdpb_inst_14.INIT_RAM_10 = 256'h9D9D9D9B9D9D9D9C9F9D9D9D9C9C9D9D9D9D9B9C9D9D9B9C9D9E9D9D9D9D9D9E;
defparam sdpb_inst_14.INIT_RAM_11 = 256'h9C9C9A9C9C9B9B9B9B9C9D9C9D9C9D9D9C9D9C9D9E9D9E9E9E9D9D9C9E9B9E9C;
defparam sdpb_inst_14.INIT_RAM_12 = 256'hA19FA0A0A0A0A0A0A0A0A0A09F9E9D9C9F9D9D9D9B9B9D9C9B9C9D9C9C9C9B9D;
defparam sdpb_inst_14.INIT_RAM_13 = 256'hA3A2A2A2A0A0A0A0A0A0A19F9FA1A0A1A1A0A09FA09FA0A09F9FA09F9FA1A0A2;
defparam sdpb_inst_14.INIT_RAM_14 = 256'h5F656D60969C9EA0A1A3A3A5A5A4A5A4A3A3A2A2A3A5A4A2A5A4A2A2A4A5A4A3;
defparam sdpb_inst_14.INIT_RAM_15 = 256'hA5A5A5A4A3A2A09F9D9C99948F8A857E70604F1049293C74CD6B5A337B787677;
defparam sdpb_inst_14.INIT_RAM_16 = 256'h9D9C9C9D9D9D9E9F9E9E9F9F9FA0A0A1A3A2A3A4A4A4A4A4A4A6A6A6A5A6A7A6;
defparam sdpb_inst_14.INIT_RAM_17 = 256'h9C9C9C9C9B9C9C9C9C9D9B9D9C9C9C9C9C9B9B9C9C9B9B9B9D9B9C9B9C9C9C9D;
defparam sdpb_inst_14.INIT_RAM_18 = 256'h9A9A9B9B9B9B9B9A9D9B9B9D9C9B9B9D9C9C9C9D9C9C9C9D9C9C9C9D9C9D9B9C;
defparam sdpb_inst_14.INIT_RAM_19 = 256'h9F9F9F9E9F9EA09FA09F9F9F9F9E9E9D9E9D9C9C9D9C9C9C9A9C9B9C9C9B9B99;
defparam sdpb_inst_14.INIT_RAM_1A = 256'hA3A3A2A2A1A19FA19E9D9FA09F9EA0A09DA0A09E9E9E9EA0A0A09F9F9E9FA09F;
defparam sdpb_inst_14.INIT_RAM_1B = 256'h6E77664C60939D9FA0A1A2A3A3A3A4A3A4A4A3A4A3A4A4A5A2A3A4A3A3A3A2A2;
defparam sdpb_inst_14.INIT_RAM_1C = 256'hA6A6A7A6A5A5A5A3A2A2A09F9D9B9894918D827C6F64544D45406881858C5F0F;
defparam sdpb_inst_14.INIT_RAM_1D = 256'h9A9C9C9B9C9C9B9D9D9D9C9D9F9EA09FA19FA0A2A2A2A3A4A4A4A4A5A6A6A6A6;
defparam sdpb_inst_14.INIT_RAM_1E = 256'h9A9A9C9B9B9B9C9B9B9C9B9A9A9A9B9B9A9A9B9B9A989A9A9C9A9A9A9A9A9B9B;
defparam sdpb_inst_14.INIT_RAM_1F = 256'h9A9A9A9B999B9A9A9A999B999A9A9A9B9B9B9B9B9A9B9B9A9B9C9B9B9B9B9B9B;
defparam sdpb_inst_14.INIT_RAM_20 = 256'h9E9C9E9E9E9E9E9F9E9F9F9F9F9F9E9F9D9D9C9B9C9C9A9C9B9A9B9A9A9C999B;
defparam sdpb_inst_14.INIT_RAM_21 = 256'hA1A1A3A1A3A09EA09F9E9D9E9D9E9D9F9E9E9E9F9E9E9F9E9EA09E9E9F9EA09E;
defparam sdpb_inst_14.INIT_RAM_22 = 256'h7C7460366161949A9DA0A3A2A3A2A3A4A5A3A3A4A3A3A4A4A3A3A1A3A3A3A3A3;
defparam sdpb_inst_14.INIT_RAM_23 = 256'hA5A5A6A5A6A5A6A6A5A5A4A4A3A29F9F9E9D9997948B847B736A63636B6E7072;
defparam sdpb_inst_14.INIT_RAM_24 = 256'h99989A9B999B9B9A9B9B9D9C9C9C9D9D9E9FA0A0A1A1A0A2A2A2A3A3A3A5A4A6;
defparam sdpb_inst_14.INIT_RAM_25 = 256'h999A9B9B9A9A999A9A9B9A989A999A9A999A9A9A9B9999999999999A999A999A;
defparam sdpb_inst_14.INIT_RAM_26 = 256'h99999A9998989999999897999A98989B99999A989A9A999B9A9A9A9B9B9A9C9A;
defparam sdpb_inst_14.INIT_RAM_27 = 256'h9D9E9D9D9C9D9D9E9D9D9E9E9D9E9E9F9D9C9E9D9C9B999B9A99989A999A9999;
defparam sdpb_inst_14.INIT_RAM_28 = 256'hA2A3A09FA1A0A2A09D9DA09E9D9E9F9E9F9D9F9D9F9D9F9D9E9D9D9D9D9C9D9D;
defparam sdpb_inst_14.INIT_RAM_29 = 256'h7072767E828C8E97999C9FA1A0A2A3A4A3A5A4A5A4A4A4A2A2A1A2A1A3A1A2A0;
defparam sdpb_inst_14.INIT_RAM_2A = 256'hA5A4A5A6A6A6A6A6A4A5A6A5A6A5A4A4A2A2A0A09E9C9B9994908E88837F7572;
defparam sdpb_inst_14.INIT_RAM_2B = 256'h9A999998989A9A989A9A9A999B999B9B9B9D9D9D9F9FA0A09FA1A1A2A2A2A3A4;
defparam sdpb_inst_14.INIT_RAM_2C = 256'h99999899989997999A989998989A9999989A9B9998999A999797989998979798;
defparam sdpb_inst_14.INIT_RAM_2D = 256'h99999998999A98969798989798969998999898999A9897999999999B9A9A9998;
defparam sdpb_inst_14.INIT_RAM_2E = 256'h9D9C9C9B9B9B9C9B9B9B9A9D9C9B9C9C9B9D9C9B999899989A99999A979A9997;
defparam sdpb_inst_14.INIT_RAM_2F = 256'hA3A0A1A0A1A0A0A09F9FA09E9C9E9E9C9C9B9B9E9D9D9C9D9B9C9C9D9C9D9A9C;
defparam sdpb_inst_14.INIT_RAM_30 = 256'h908E8C8B8E8F9295989A9DA0A0A3A2A1A3A4A4A3A3A3A2A2A3A2A1A2A2A2A1A1;
defparam sdpb_inst_14.INIT_RAM_31 = 256'hA2A3A3A3A4A4A5A4A5A6A6A6A5A5A7A5A3A5A5A4A4A3A2A09F9E9C9B98969492;
defparam sdpb_inst_14.INIT_RAM_32 = 256'h97969795999797979798999899999A9B9B999B9C9C9C9D9E9EA0A0A1A0A0A1A1;
defparam sdpb_inst_14.INIT_RAM_33 = 256'h9897989799979997999998989798989999999798989798979897989897979698;
defparam sdpb_inst_14.INIT_RAM_34 = 256'h9996989896969897989895969799969796969798979797989997999899979999;
defparam sdpb_inst_14.INIT_RAM_35 = 256'h9C9B9C9C9B9B9B9B999A9A9B9D9B9C9B9A9B9B9B989998989797979898989897;
defparam sdpb_inst_14.INIT_RAM_36 = 256'hA2A2A2A1A1A0A2A1A09FA19D9F9D9C9D9E9A9B9A9A9C9C9C9D9B9D9E9B9C9B9D;
defparam sdpb_inst_14.INIT_RAM_37 = 256'h9B9A9B97989A96989A9C9C9EA0A09EA2A4A4A3A4A5A4A2A2A2A1A3A2A3A29FA0;
defparam sdpb_inst_14.INIT_RAM_38 = 256'hA1A1A2A3A1A3A3A4A4A6A4A6A4A5A6A6A5A5A6A5A5A4A4A4A4A3A4A2A09E9D9D;
defparam sdpb_inst_14.INIT_RAM_39 = 256'h959596969396979495969797979797999A999A9A99999C9B9B9C9D9E9DA09EA0;
defparam sdpb_inst_14.INIT_RAM_3A = 256'h9996989697969796969796989798979597979599969594959797969595959796;
defparam sdpb_inst_14.INIT_RAM_3B = 256'h9495959697949597989895969797959797969796969797979897959698989497;
defparam sdpb_inst_14.INIT_RAM_3C = 256'h9A9C9B9A9A9A979999999B999A999A989A989896999898969898979596959596;
defparam sdpb_inst_14.INIT_RAM_3D = 256'h000000000000000000000000000000000000009A9B999A9B989C9D9A9D999C99;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clkb),
  .CE(oce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[13]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clkb),
  .CE(oce)
);
DFFE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb)
);
DFFE dff_inst_5 (
  .Q(dff_q_5),
  .D(dff_q_4),
  .CLK(clkb),
  .CE(oce)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(sdpb_inst_12_dout[0]),
  .I1(sdpb_inst_14_dout[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(sdpb_inst_8_dout[0]),
  .I1(mux_o_6),
  .S0(dff_q_3)
);
MUX2 mux_inst_9 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(mux_o_8),
  .S0(dff_q_1)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(sdpb_inst_12_dout[1]),
  .I1(sdpb_inst_14_dout[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(sdpb_inst_8_dout[1]),
  .I1(mux_o_16),
  .S0(dff_q_3)
);
MUX2 mux_inst_19 (
  .O(dout[1]),
  .I0(sdpb_inst_1_dout[1]),
  .I1(mux_o_18),
  .S0(dff_q_1)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(sdpb_inst_12_dout[2]),
  .I1(sdpb_inst_14_dout[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(sdpb_inst_9_dout[2]),
  .I1(mux_o_26),
  .S0(dff_q_3)
);
MUX2 mux_inst_29 (
  .O(dout[2]),
  .I0(sdpb_inst_2_dout[2]),
  .I1(mux_o_28),
  .S0(dff_q_1)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(sdpb_inst_12_dout[3]),
  .I1(sdpb_inst_14_dout[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(sdpb_inst_9_dout[3]),
  .I1(mux_o_36),
  .S0(dff_q_3)
);
MUX2 mux_inst_39 (
  .O(dout[3]),
  .I0(sdpb_inst_3_dout[3]),
  .I1(mux_o_38),
  .S0(dff_q_1)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sdpb_inst_13_dout[4]),
  .I1(sdpb_inst_14_dout[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(sdpb_inst_10_dout[4]),
  .I1(mux_o_46),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(dout[4]),
  .I0(sdpb_inst_4_dout[4]),
  .I1(mux_o_48),
  .S0(dff_q_1)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(sdpb_inst_13_dout[5]),
  .I1(sdpb_inst_14_dout[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(sdpb_inst_10_dout[5]),
  .I1(mux_o_56),
  .S0(dff_q_3)
);
MUX2 mux_inst_59 (
  .O(dout[5]),
  .I0(sdpb_inst_5_dout[5]),
  .I1(mux_o_58),
  .S0(dff_q_1)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(sdpb_inst_13_dout[6]),
  .I1(sdpb_inst_14_dout[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(sdpb_inst_11_dout[6]),
  .I1(mux_o_66),
  .S0(dff_q_3)
);
MUX2 mux_inst_69 (
  .O(dout[6]),
  .I0(sdpb_inst_6_dout[6]),
  .I1(mux_o_68),
  .S0(dff_q_1)
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(sdpb_inst_13_dout[7]),
  .I1(sdpb_inst_14_dout[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(sdpb_inst_11_dout[7]),
  .I1(mux_o_76),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(dout[7]),
  .I0(sdpb_inst_7_dout[7]),
  .I1(mux_o_78),
  .S0(dff_q_1)
);
endmodule //Gowin_SDPB5
